------------------------------------------------------------------------------
--  This file is a part of the GRLIB VHDL IP LIBRARY
--  Copyright (C) 2009, Aeroflex Gaisler AB - all rights reserved.
--
-- ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN 
-- ACCORDANCE WITH THE GAISLER LICENSE AGREEMENT AND MUST BE APPROVED 
-- IN ADVANCE IN WRITING.
------------------------------------------------------------------------------
--
-- Written by Synplicity
-- Product Version "E-2010.09"
-- Program "Synplify Pro", Mapper "maprc, Build 140R"
-- Mon Jan 31 16:12:40 2011
--

--
-- Written by Synplify Pro version Build 140R
-- Mon Jan 31 16:12:40 2011
--

--
library ieee, stratixiii;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
--library synplify;
--use synplify.components.all;
use stratixiii.stratixiii_components.all;
library altera;
use altera.altera_primitives_components.all;

entity grlfpw_0_stratixiii is
port(
  rst :  in std_logic;
  clk :  in std_logic;
  holdn :  in std_logic;
  cpi_flush :  in std_logic;
  cpi_exack :  in std_logic;
  cpi_a_rs1 : in std_logic_vector(4 downto 0);
  cpi_d_pc : in std_logic_vector(31 downto 0);
  cpi_d_inst : in std_logic_vector(31 downto 0);
  cpi_d_cnt : in std_logic_vector(1 downto 0);
  cpi_d_trap :  in std_logic;
  cpi_d_annul :  in std_logic;
  cpi_d_pv :  in std_logic;
  cpi_a_pc : in std_logic_vector(31 downto 0);
  cpi_a_inst : in std_logic_vector(31 downto 0);
  cpi_a_cnt : in std_logic_vector(1 downto 0);
  cpi_a_trap :  in std_logic;
  cpi_a_annul :  in std_logic;
  cpi_a_pv :  in std_logic;
  cpi_e_pc : in std_logic_vector(31 downto 0);
  cpi_e_inst : in std_logic_vector(31 downto 0);
  cpi_e_cnt : in std_logic_vector(1 downto 0);
  cpi_e_trap :  in std_logic;
  cpi_e_annul :  in std_logic;
  cpi_e_pv :  in std_logic;
  cpi_m_pc : in std_logic_vector(31 downto 0);
  cpi_m_inst : in std_logic_vector(31 downto 0);
  cpi_m_cnt : in std_logic_vector(1 downto 0);
  cpi_m_trap :  in std_logic;
  cpi_m_annul :  in std_logic;
  cpi_m_pv :  in std_logic;
  cpi_x_pc : in std_logic_vector(31 downto 0);
  cpi_x_inst : in std_logic_vector(31 downto 0);
  cpi_x_cnt : in std_logic_vector(1 downto 0);
  cpi_x_trap :  in std_logic;
  cpi_x_annul :  in std_logic;
  cpi_x_pv :  in std_logic;
  cpi_lddata : in std_logic_vector(31 downto 0);
  cpi_dbg_enable :  in std_logic;
  cpi_dbg_write :  in std_logic;
  cpi_dbg_fsr :  in std_logic;
  cpi_dbg_addr : in std_logic_vector(4 downto 0);
  cpi_dbg_data : in std_logic_vector(31 downto 0);
  cpo_data : out std_logic_vector(31 downto 0);
  cpo_exc :  out std_logic;
  cpo_cc : out std_logic_vector(1 downto 0);
  cpo_ccv :  out std_logic;
  cpo_ldlock :  out std_logic;
  cpo_holdn :  out std_logic;
  cpo_dbg_data : out std_logic_vector(31 downto 0);
  rfi1_rd1addr : out std_logic_vector(3 downto 0);
  rfi1_rd2addr : out std_logic_vector(3 downto 0);
  rfi1_wraddr : out std_logic_vector(3 downto 0);
  rfi1_wrdata : out std_logic_vector(31 downto 0);
  rfi1_ren1 :  out std_logic;
  rfi1_ren2 :  out std_logic;
  rfi1_wren :  out std_logic;
  rfi2_rd1addr : out std_logic_vector(3 downto 0);
  rfi2_rd2addr : out std_logic_vector(3 downto 0);
  rfi2_wraddr : out std_logic_vector(3 downto 0);
  rfi2_wrdata : out std_logic_vector(31 downto 0);
  rfi2_ren1 :  out std_logic;
  rfi2_ren2 :  out std_logic;
  rfi2_wren :  out std_logic;
  rfo1_data1 : in std_logic_vector(31 downto 0);
  rfo1_data2 : in std_logic_vector(31 downto 0);
  rfo2_data1 : in std_logic_vector(31 downto 0);
  rfo2_data2 : in std_logic_vector(31 downto 0));
end grlfpw_0_stratixiii;

architecture beh of grlfpw_0_stratixiii is
  signal devclrn : std_logic := '1';
  signal devpor : std_logic := '1';
  signal devoe : std_logic := '0';
  signal \GRLFPC2_0.FPI.OP2\ : std_logic_vector(63 downto 32);
  signal \GRLFPC2_0.R.FSR.RD\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.FPO.FRAC\ : std_logic_vector(54 downto 3);
  signal \GRLFPC2_0.FPO.EXP\ : std_logic_vector(10 downto 0);
  signal \GRLFPC2_0.R.STATE\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.R.I.INST\ : std_logic_vector(31 downto 0);
  signal \GRLFPC2_0.R.FSR.TEM\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.R.I.EXC\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.R.FSR.AEXC\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.R.A.RS1\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.R.A.RS2\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.R.FSR.CEXC\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.R.FSR.FTT\ : std_logic_vector(2 downto 0);
  signal \GRLFPC2_0.R.I.RES\ : std_logic_vector(63 downto 0);
  signal \GRLFPC2_0.COMB.V.I.RES_1\ : std_logic_vector(63 to 63);
  signal \GRLFPC2_0.R.A.RF1REN\ : std_logic_vector(2 downto 1);
  signal \GRLFPC2_0.R.A.RF2REN\ : std_logic_vector(2 downto 1);
  signal \GRLFPC2_0.R.I.CC\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.FPCI_O\ : std_logic_vector(314 downto 0);
  signal \GRLFPC2_0.R.STATE_O\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.FPCI_O_3\ : std_logic_vector(74 downto 0);
  signal \GRLFPC2_0.R.STATE_O_3\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.FPCI_O_0\ : std_logic_vector(70 downto 59);
  signal \GRLFPC2_0.R.I.PC_O\ : std_logic_vector(31 downto 2);
  signal \GRLFPC2_0.R.I.EXC_MB\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.COMB.RS1_1\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.COMB.RS2_1\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\ : std_logic_vector(85 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\ : std_logic_vector(16 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\ : std_logic_vector(377 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\ : std_logic_vector(57 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\ : std_logic_vector(57 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\ : std_logic_vector(12 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_57\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_56\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_55\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_54\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_53\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_52\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_51\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_50\ : std_logic_vector(7 to 7);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_49\ : std_logic_vector(8 to 8);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_48\ : std_logic_vector(9 to 9);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_47\ : std_logic_vector(10 to 10);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_46\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_45\ : std_logic_vector(12 to 12);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_44\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_43\ : std_logic_vector(14 to 14);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_42\ : std_logic_vector(15 to 15);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_41\ : std_logic_vector(16 to 16);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_40\ : std_logic_vector(17 to 17);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_39\ : std_logic_vector(18 to 18);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_38\ : std_logic_vector(19 to 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_37\ : std_logic_vector(20 to 20);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_36\ : std_logic_vector(21 to 21);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_35\ : std_logic_vector(22 to 22);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_34\ : std_logic_vector(23 to 23);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_33\ : std_logic_vector(24 to 24);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_32\ : std_logic_vector(25 to 25);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_31\ : std_logic_vector(26 to 26);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_30\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_29\ : std_logic_vector(28 to 28);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_28\ : std_logic_vector(29 to 29);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_27\ : std_logic_vector(30 to 30);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_26\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_25\ : std_logic_vector(32 to 32);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_24\ : std_logic_vector(33 to 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_23\ : std_logic_vector(34 to 34);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_22\ : std_logic_vector(35 to 35);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_21\ : std_logic_vector(36 to 36);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_20\ : std_logic_vector(37 to 37);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_19\ : std_logic_vector(38 to 38);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_18\ : std_logic_vector(39 to 39);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_17\ : std_logic_vector(40 to 40);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_16\ : std_logic_vector(41 to 41);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_15\ : std_logic_vector(42 to 42);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_14\ : std_logic_vector(43 to 43);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_13\ : std_logic_vector(44 to 44);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_12\ : std_logic_vector(45 to 45);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_11\ : std_logic_vector(46 to 46);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_10\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_9\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_8\ : std_logic_vector(49 to 49);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_7\ : std_logic_vector(50 to 50);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_6\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_5\ : std_logic_vector(52 to 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_113\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SBLSBS_1\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_112\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_111\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_110\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_109\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_108\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_107\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_106\ : std_logic_vector(7 to 7);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_105\ : std_logic_vector(8 to 8);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_104\ : std_logic_vector(9 to 9);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_103\ : std_logic_vector(10 to 10);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_102\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_101\ : std_logic_vector(12 to 12);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_100\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_99\ : std_logic_vector(14 to 14);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_98\ : std_logic_vector(15 to 15);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_97\ : std_logic_vector(16 to 16);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_96\ : std_logic_vector(17 to 17);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_95\ : std_logic_vector(18 to 18);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_94\ : std_logic_vector(19 to 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_93\ : std_logic_vector(20 to 20);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_92\ : std_logic_vector(21 to 21);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_91\ : std_logic_vector(22 to 22);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_90\ : std_logic_vector(23 to 23);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_89\ : std_logic_vector(24 to 24);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_88\ : std_logic_vector(25 to 25);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_87\ : std_logic_vector(26 to 26);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_86\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_85\ : std_logic_vector(28 to 28);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_84\ : std_logic_vector(29 to 29);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_83\ : std_logic_vector(30 to 30);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_82\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_81\ : std_logic_vector(32 to 32);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_80\ : std_logic_vector(33 to 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_79\ : std_logic_vector(34 to 34);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_78\ : std_logic_vector(35 to 35);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_77\ : std_logic_vector(36 to 36);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_76\ : std_logic_vector(37 to 37);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_75\ : std_logic_vector(38 to 38);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_74\ : std_logic_vector(39 to 39);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_73\ : std_logic_vector(40 to 40);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_72\ : std_logic_vector(41 to 41);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_71\ : std_logic_vector(42 to 42);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_70\ : std_logic_vector(43 to 43);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_69\ : std_logic_vector(44 to 44);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_68\ : std_logic_vector(45 to 45);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_67\ : std_logic_vector(46 to 46);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_66\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_65\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_64\ : std_logic_vector(49 to 49);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_63\ : std_logic_vector(50 to 50);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_62\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\ : std_logic_vector(57 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SCLSBS_2\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SCLSBS_1\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_168\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_167\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_166\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_165\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_164\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_163\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_162\ : std_logic_vector(7 to 7);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_161\ : std_logic_vector(8 to 8);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_160\ : std_logic_vector(9 to 9);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_159\ : std_logic_vector(10 to 10);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_158\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_157\ : std_logic_vector(12 to 12);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_156\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_155\ : std_logic_vector(14 to 14);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_154\ : std_logic_vector(15 to 15);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_153\ : std_logic_vector(16 to 16);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_152\ : std_logic_vector(17 to 17);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_151\ : std_logic_vector(18 to 18);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_150\ : std_logic_vector(19 to 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_149\ : std_logic_vector(20 to 20);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_148\ : std_logic_vector(21 to 21);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_147\ : std_logic_vector(22 to 22);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_146\ : std_logic_vector(23 to 23);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_145\ : std_logic_vector(24 to 24);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_144\ : std_logic_vector(25 to 25);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_143\ : std_logic_vector(26 to 26);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_142\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_141\ : std_logic_vector(28 to 28);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_140\ : std_logic_vector(29 to 29);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_139\ : std_logic_vector(30 to 30);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_138\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_137\ : std_logic_vector(32 to 32);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_136\ : std_logic_vector(33 to 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_135\ : std_logic_vector(34 to 34);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_134\ : std_logic_vector(35 to 35);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_133\ : std_logic_vector(36 to 36);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_132\ : std_logic_vector(37 to 37);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_131\ : std_logic_vector(38 to 38);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_130\ : std_logic_vector(39 to 39);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_129\ : std_logic_vector(40 to 40);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_128\ : std_logic_vector(41 to 41);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_127\ : std_logic_vector(42 to 42);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_126\ : std_logic_vector(43 to 43);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_125\ : std_logic_vector(44 to 44);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_124\ : std_logic_vector(45 to 45);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_123\ : std_logic_vector(46 to 46);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_122\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_121\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_120\ : std_logic_vector(49 to 49);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_119\ : std_logic_vector(50 to 50);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW_2\ : std_logic_vector(65 to 65);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\ : std_logic_vector(55 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\ : std_logic_vector(112 downto 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\ : std_logic_vector(9 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\ : std_logic_vector(2 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\ : std_logic_vector(12 downto 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_DIVMULTV\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\ : std_logic_vector(375 downto 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_14\ : std_logic_vector(172 downto 141);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\ : std_logic_vector(83 downto 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SCTRL_NEW\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW_6\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\ : std_logic_vector(112 downto 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19\ : std_logic_vector(9 to 9);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.CONDITIONAL\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_D\ : std_logic_vector(7 to 7);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1\ : std_logic_vector(45 to 45);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\ : std_logic_vector(113 downto 58);
  signal \GRLFPC2_0.R.I.PC\ : std_logic_vector(26 downto 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\ : std_logic_vector(56 downto 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\ : std_logic_vector(48 downto 12);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\ : std_logic_vector(57 downto 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\ : std_logic_vector(45 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\ : std_logic_vector(54 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\ : std_logic_vector(257 to 257);
  signal \GRLFPC2_0.FPI.OP1\ : std_logic_vector(62 downto 32);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\ : std_logic_vector(4 downto 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\ : std_logic_vector(8 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SBLSBS_2\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SALSBS_1\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SALSBS_2\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\ : std_logic_vector(8 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\ : std_logic_vector(9 downto 2);
  signal \GRLFPC2_0.COMB.V.A.RF1REN_1\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.COMB.V.A.RF2REN_1\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.COMB.WRDATA_4\ : std_logic_vector(62 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\ : std_logic_vector(115 downto 71);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\ : std_logic_vector(115 downto 71);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\ : std_logic_vector(21 downto 16);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\ : std_logic_vector(51 downto 46);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\ : std_logic_vector(6 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8_0\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_116\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_I_M\ : std_logic_vector(12 to 12);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_60\ : std_logic_vector(53 to 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A32_18_1\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_32_1\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_12\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_8\ : std_logic_vector(60 downto 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_A2_14_S\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_A2_5_S\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_A2_3_S\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_10_TZ\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_IV_1_TZ\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_A2_2_3\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_1_TZ\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_3_0\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_13_1\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_15_1\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A32_19_0\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_6_1\ : std_logic_vector(59 downto 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_4_1\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_32_1\ : std_logic_vector(58 to 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7_0\ : std_logic_vector(52 to 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_16_0\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A32_1_0\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A8_2_0\ : std_logic_vector(62 to 62);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_I_I_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_3_I\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\ : std_logic_vector(56 downto 9);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\ : std_logic_vector(55 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\ : std_logic_vector(45 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\ : std_logic_vector(55 downto 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_I_O2_3_0\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_O2_10_4\ : std_logic_vector(83 to 83);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_I_O2_4_4\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_O2_12_4\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_O2_11_3\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_6_1_0\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_7_1\ : std_logic_vector(53 to 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A32_13_1_0\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_1_1\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_15_0\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_15_0\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A32_3_1\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A32_2_0\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_37_0\ : std_logic_vector(19 to 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_4_1\ : std_logic_vector(33 to 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11_1\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_28_0\ : std_logic_vector(19 to 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_23_0\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_5_0\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_26_0\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_8_0\ : std_logic_vector(18 to 18);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_11_0\ : std_logic_vector(32 to 32);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A8_5_0\ : std_logic_vector(62 to 62);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A11_3_0\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A11_3_1\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_28_0\ : std_logic_vector(58 to 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_28_1\ : std_logic_vector(58 to 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_4_1\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_0_1\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_10_0\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_0_0\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_52_0\ : std_logic_vector(58 to 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_52_1\ : std_logic_vector(58 to 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_1\ : std_logic_vector(26 to 26);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A11_5_2\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A11_5_3\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_33_0\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A32_11_0\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A28_0_1\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7_3_0\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A28_4_1\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_3_1\ : std_logic_vector(25 to 25);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_3_0\ : std_logic_vector(52 to 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A28_8_0\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_1_1\ : std_logic_vector(33 to 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_2_0_0\ : std_logic_vector(36 to 36);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_A28_6_0\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_13_0\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_9_0_0\ : std_logic_vector(53 to 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_3_1\ : std_logic_vector(32 to 32);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_2_1\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A26_12_0\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A28_7_0\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_27_0\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_A28_5_1\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_4_0\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_3_0\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_8_0\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_8_1\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A32_8_0\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A32_0\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_34_0\ : std_logic_vector(58 to 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_26_1\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_0_0\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_2_0\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_I_O2_0\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\ : std_logic_vector(7 downto 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_5_1\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_1_2\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0_1\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A21_0\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_11_0\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1_A2_0\ : std_logic_vector(39 to 39);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A9_4_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_4_0\ : std_logic_vector(12 to 12);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_1_0\ : std_logic_vector(53 to 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0_1\ : std_logic_vector(37 to 37);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A24_0\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0_0\ : std_logic_vector(10 to 10);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_0_0\ : std_logic_vector(39 to 39);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_0\ : std_logic_vector(8 to 8);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_0\ : std_logic_vector(60 downto 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_1\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_2\ : std_logic_vector(60 downto 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_7\ : std_logic_vector(47 downto 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_9\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_11\ : std_logic_vector(60 downto 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_14\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_18\ : std_logic_vector(60 downto 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_20\ : std_logic_vector(60 downto 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_22\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_3\ : std_logic_vector(60 downto 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_6\ : std_logic_vector(60 downto 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_13\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_16\ : std_logic_vector(60 downto 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_17\ : std_logic_vector(60 downto 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_21\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_4\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_5\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_19\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_A2_7_1\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_1\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV_0\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_A2_41_0\ : std_logic_vector(83 to 83);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_A2_41_2\ : std_logic_vector(83 to 83);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_O2_4_0\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_A2_7_0\ : std_logic_vector(83 to 83);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_A2_7_2\ : std_logic_vector(83 to 83);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_0\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0\ : std_logic_vector(9 to 9);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0_0\ : std_logic_vector(7 to 7);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_A2_1_A2_2\ : std_logic_vector(83 to 83);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_A2_1_A2_7\ : std_logic_vector(83 to 83);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_A2_1_A2_9\ : std_logic_vector(83 to 83);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8_I\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.EXTEND.TEMP_0\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\ : std_logic_vector(30 downto 9);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\ : std_logic_vector(85 downto 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO\ : std_logic_vector(7 downto 0);
  signal CPI_D_INST_RETO : std_logic_vector(12 downto 5);
  signal RFO2_DATA1_RETO : std_logic_vector(28 downto 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\ : std_logic_vector(109 downto 64);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5_RETI\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M11\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1_RETO\ : std_logic_vector(115 downto 71);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0_RETO\ : std_logic_vector(115 downto 71);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_3_I_RETO\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.FPO.FRAC_RETO\ : std_logic_vector(5 downto 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\ : std_logic_vector(51 downto 50);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\ : std_logic_vector(113 downto 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_I_O2_4_4_RETI\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2_RETI\ : std_logic_vector(9 to 9);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\ : std_logic_vector(80 downto 64);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\ : std_logic_vector(72 downto 71);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW\ : std_logic_vector(7 to 7);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\ : std_logic_vector(65 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\ : std_logic_vector(65 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\ : std_logic_vector(43 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\ : std_logic_vector(42 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\ : std_logic_vector(42 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI_0\ : std_logic_vector(10 to 10);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\ : std_logic_vector(84 downto 78);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\ : std_logic_vector(81 downto 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\ : std_logic_vector(244 downto 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\ : std_logic_vector(3 downto 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\ : std_logic_vector(243 downto 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_0\ : std_logic_vector(15 to 15);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\ : std_logic_vector(3 downto 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_1\ : std_logic_vector(15 to 15);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_2\ : std_logic_vector(15 to 15);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_3\ : std_logic_vector(15 to 15);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_4\ : std_logic_vector(15 to 15);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\ : std_logic_vector(42 downto 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_5\ : std_logic_vector(15 to 15);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\ : std_logic_vector(8 downto 2);
  signal \GRLFPC2_0.R.STATE_O_3_0\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\ : std_logic_vector(8 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\ : std_logic_vector(57 downto 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_0\ : std_logic_vector(7 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_3\ : std_logic_vector(57 downto 23);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_1\ : std_logic_vector(5 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_4\ : std_logic_vector(55 downto 23);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_6\ : std_logic_vector(42 downto 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_6\ : std_logic_vector(15 to 15);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\ : std_logic_vector(84 downto 78);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO_0\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO_0\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_0\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\ : std_logic_vector(84 downto 78);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO_1\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO_1\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_1\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\ : std_logic_vector(84 downto 78);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO_2\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO_2\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_2\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\ : std_logic_vector(84 downto 78);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO_3\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO_3\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_3\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\ : std_logic_vector(84 downto 78);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO_4\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO_4\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_4\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO_5\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO_5\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_5\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\ : std_logic_vector(84 downto 83);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO_6\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO_6\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_6\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\ : std_logic_vector(84 downto 83);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO_7\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO_7\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_7\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\ : std_logic_vector(81 to 81);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\ : std_logic_vector(84 downto 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\ : std_logic_vector(81 to 81);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\ : std_logic_vector(84 downto 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\ : std_logic_vector(81 to 81);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_2\ : std_logic_vector(84 downto 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_3\ : std_logic_vector(84 downto 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\ : std_logic_vector(81 downto 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_4\ : std_logic_vector(84 downto 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\ : std_logic_vector(81 downto 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_5\ : std_logic_vector(84 downto 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\ : std_logic_vector(81 downto 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_6\ : std_logic_vector(84 downto 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\ : std_logic_vector(81 downto 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_7\ : std_logic_vector(84 downto 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\ : std_logic_vector(81 downto 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_8\ : std_logic_vector(84 downto 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\ : std_logic_vector(85 downto 83);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_0\ : std_logic_vector(7 downto 0);
  signal CPI_D_INST_RETO_0 : std_logic_vector(12 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\ : std_logic_vector(85 downto 83);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_1\ : std_logic_vector(7 downto 0);
  signal CPI_D_INST_RETO_1 : std_logic_vector(12 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\ : std_logic_vector(85 downto 83);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_2\ : std_logic_vector(7 downto 0);
  signal CPI_D_INST_RETO_2 : std_logic_vector(12 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\ : std_logic_vector(85 to 85);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_3\ : std_logic_vector(7 downto 0);
  signal CPI_D_INST_RETO_3 : std_logic_vector(12 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\ : std_logic_vector(85 to 85);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_4\ : std_logic_vector(7 downto 0);
  signal CPI_D_INST_RETO_4 : std_logic_vector(12 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\ : std_logic_vector(85 to 85);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_5\ : std_logic_vector(7 downto 0);
  signal CPI_D_INST_RETO_5 : std_logic_vector(12 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\ : std_logic_vector(85 to 85);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_6\ : std_logic_vector(7 downto 0);
  signal CPI_D_INST_RETO_6 : std_logic_vector(12 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\ : std_logic_vector(85 to 85);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_7\ : std_logic_vector(7 downto 0);
  signal CPI_D_INST_RETO_7 : std_logic_vector(12 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\ : std_logic_vector(85 to 85);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_8\ : std_logic_vector(7 downto 0);
  signal CPI_D_INST_RETO_8 : std_logic_vector(12 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\ : std_logic_vector(80 downto 78);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\ : std_logic_vector(80 downto 78);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\ : std_logic_vector(80 downto 78);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_9\ : std_logic_vector(3 downto 0);
  signal CPI_D_INST_RETO_9 : std_logic_vector(11 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_9\ : std_logic_vector(79 to 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_10\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_10\ : std_logic_vector(79 to 79);
  signal CPI_D_INST_RETO_10 : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\ : std_logic_vector(83 to 83);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\ : std_logic_vector(83 to 83);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\ : std_logic_vector(83 to 83);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\ : std_logic_vector(82 to 82);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_0\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\ : std_logic_vector(82 to 82);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_1\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\ : std_logic_vector(82 to 82);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_2\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\ : std_logic_vector(82 to 82);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_3\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\ : std_logic_vector(82 to 82);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_4\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\ : std_logic_vector(82 to 82);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_5\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\ : std_logic_vector(82 to 82);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_6\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\ : std_logic_vector(82 to 82);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_7\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\ : std_logic_vector(82 to 82);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_8\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\ : std_logic_vector(82 to 82);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_9\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_5\ : std_logic_vector(55 downto 23);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260_0\ : std_logic_vector(84 to 84);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272_0\ : std_logic_vector(85 to 85);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_7\ : std_logic_vector(42 to 42);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_7\ : std_logic_vector(15 to 15);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_2\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_3\ : std_logic_vector(4 to 4);
  signal CPO_DATAZ : std_logic_vector(31 downto 0);
  signal CPO_CCZ : std_logic_vector(1 downto 0);
  signal CPO_DBG_DATAZ : std_logic_vector(31 downto 0);
  signal RFI1_WRDATAZ : std_logic_vector(31 downto 0);
  signal RFI2_RD1ADDRZ : std_logic_vector(3 downto 0);
  signal RFI2_RD2ADDRZ : std_logic_vector(3 downto 0);
  signal RFI2_WRADDRZ : std_logic_vector(3 downto 0);
  signal RFI2_WRDATAZ : std_logic_vector(31 downto 0);
  signal RST_INTERNAL : std_logic ;
  signal CLK_INTERNAL : std_logic ;
  signal HOLDN_INTERNAL : std_logic ;
  signal CPI_FLUSH_INTERNAL : std_logic ;
  signal CPI_EXACK_INTERNAL : std_logic ;
  signal CPI_A_RS1_INTERNAL : std_logic ;
  signal CPI_A_RS1_INTERNAL_0 : std_logic ;
  signal CPI_A_RS1_INTERNAL_1 : std_logic ;
  signal CPI_A_RS1_INTERNAL_2 : std_logic ;
  signal CPI_A_RS1_INTERNAL_3 : std_logic ;
  signal CPI_D_PC_INTERNAL : std_logic ;
  signal CPI_D_PC_INTERNAL_0 : std_logic ;
  signal CPI_D_PC_INTERNAL_1 : std_logic ;
  signal CPI_D_PC_INTERNAL_2 : std_logic ;
  signal CPI_D_PC_INTERNAL_3 : std_logic ;
  signal CPI_D_PC_INTERNAL_4 : std_logic ;
  signal CPI_D_PC_INTERNAL_5 : std_logic ;
  signal CPI_D_PC_INTERNAL_6 : std_logic ;
  signal CPI_D_PC_INTERNAL_7 : std_logic ;
  signal CPI_D_PC_INTERNAL_8 : std_logic ;
  signal CPI_D_PC_INTERNAL_9 : std_logic ;
  signal CPI_D_PC_INTERNAL_10 : std_logic ;
  signal CPI_D_PC_INTERNAL_11 : std_logic ;
  signal CPI_D_PC_INTERNAL_12 : std_logic ;
  signal CPI_D_PC_INTERNAL_13 : std_logic ;
  signal CPI_D_PC_INTERNAL_14 : std_logic ;
  signal CPI_D_PC_INTERNAL_15 : std_logic ;
  signal CPI_D_PC_INTERNAL_16 : std_logic ;
  signal CPI_D_PC_INTERNAL_17 : std_logic ;
  signal CPI_D_PC_INTERNAL_18 : std_logic ;
  signal CPI_D_PC_INTERNAL_19 : std_logic ;
  signal CPI_D_PC_INTERNAL_20 : std_logic ;
  signal CPI_D_PC_INTERNAL_21 : std_logic ;
  signal CPI_D_PC_INTERNAL_22 : std_logic ;
  signal CPI_D_PC_INTERNAL_23 : std_logic ;
  signal CPI_D_PC_INTERNAL_24 : std_logic ;
  signal CPI_D_PC_INTERNAL_25 : std_logic ;
  signal CPI_D_PC_INTERNAL_26 : std_logic ;
  signal CPI_D_PC_INTERNAL_27 : std_logic ;
  signal CPI_D_PC_INTERNAL_28 : std_logic ;
  signal CPI_D_PC_INTERNAL_29 : std_logic ;
  signal CPI_D_PC_INTERNAL_30 : std_logic ;
  signal CPI_D_INST_INTERNAL : std_logic ;
  signal CPI_D_INST_INTERNAL_0 : std_logic ;
  signal CPI_D_INST_INTERNAL_1 : std_logic ;
  signal CPI_D_INST_INTERNAL_2 : std_logic ;
  signal CPI_D_INST_INTERNAL_3 : std_logic ;
  signal CPI_D_INST_INTERNAL_4 : std_logic ;
  signal CPI_D_INST_INTERNAL_5 : std_logic ;
  signal CPI_D_INST_INTERNAL_7 : std_logic ;
  signal CPI_D_INST_INTERNAL_8 : std_logic ;
  signal CPI_D_INST_INTERNAL_9 : std_logic ;
  signal CPI_D_INST_INTERNAL_10 : std_logic ;
  signal CPI_D_INST_INTERNAL_11 : std_logic ;
  signal CPI_D_INST_INTERNAL_12 : std_logic ;
  signal CPI_D_INST_INTERNAL_13 : std_logic ;
  signal CPI_D_INST_INTERNAL_14 : std_logic ;
  signal CPI_D_INST_INTERNAL_15 : std_logic ;
  signal CPI_D_INST_INTERNAL_16 : std_logic ;
  signal CPI_D_INST_INTERNAL_17 : std_logic ;
  signal CPI_D_INST_INTERNAL_18 : std_logic ;
  signal CPI_D_INST_INTERNAL_19 : std_logic ;
  signal CPI_D_INST_INTERNAL_20 : std_logic ;
  signal CPI_D_INST_INTERNAL_21 : std_logic ;
  signal CPI_D_INST_INTERNAL_22 : std_logic ;
  signal CPI_D_INST_INTERNAL_23 : std_logic ;
  signal CPI_D_INST_INTERNAL_24 : std_logic ;
  signal CPI_D_INST_INTERNAL_25 : std_logic ;
  signal CPI_D_INST_INTERNAL_26 : std_logic ;
  signal CPI_D_INST_INTERNAL_27 : std_logic ;
  signal CPI_D_INST_INTERNAL_28 : std_logic ;
  signal CPI_D_INST_INTERNAL_29 : std_logic ;
  signal CPI_D_INST_INTERNAL_30 : std_logic ;
  signal CPI_D_CNT_INTERNAL : std_logic ;
  signal CPI_D_CNT_INTERNAL_0 : std_logic ;
  signal CPI_D_TRAP_INTERNAL : std_logic ;
  signal CPI_D_ANNUL_INTERNAL : std_logic ;
  signal CPI_D_PV_INTERNAL : std_logic ;
  signal CPI_A_PC_INTERNAL : std_logic ;
  signal CPI_A_PC_INTERNAL_0 : std_logic ;
  signal CPI_A_PC_INTERNAL_1 : std_logic ;
  signal CPI_A_PC_INTERNAL_2 : std_logic ;
  signal CPI_A_PC_INTERNAL_3 : std_logic ;
  signal CPI_A_PC_INTERNAL_4 : std_logic ;
  signal CPI_A_PC_INTERNAL_5 : std_logic ;
  signal CPI_A_PC_INTERNAL_6 : std_logic ;
  signal CPI_A_PC_INTERNAL_7 : std_logic ;
  signal CPI_A_PC_INTERNAL_8 : std_logic ;
  signal CPI_A_PC_INTERNAL_9 : std_logic ;
  signal CPI_A_PC_INTERNAL_10 : std_logic ;
  signal CPI_A_PC_INTERNAL_11 : std_logic ;
  signal CPI_A_PC_INTERNAL_12 : std_logic ;
  signal CPI_A_PC_INTERNAL_13 : std_logic ;
  signal CPI_A_PC_INTERNAL_14 : std_logic ;
  signal CPI_A_PC_INTERNAL_15 : std_logic ;
  signal CPI_A_PC_INTERNAL_16 : std_logic ;
  signal CPI_A_PC_INTERNAL_17 : std_logic ;
  signal CPI_A_PC_INTERNAL_18 : std_logic ;
  signal CPI_A_PC_INTERNAL_19 : std_logic ;
  signal CPI_A_PC_INTERNAL_20 : std_logic ;
  signal CPI_A_PC_INTERNAL_21 : std_logic ;
  signal CPI_A_PC_INTERNAL_22 : std_logic ;
  signal CPI_A_PC_INTERNAL_23 : std_logic ;
  signal CPI_A_PC_INTERNAL_24 : std_logic ;
  signal CPI_A_PC_INTERNAL_25 : std_logic ;
  signal CPI_A_PC_INTERNAL_26 : std_logic ;
  signal CPI_A_PC_INTERNAL_27 : std_logic ;
  signal CPI_A_PC_INTERNAL_28 : std_logic ;
  signal CPI_A_PC_INTERNAL_29 : std_logic ;
  signal CPI_A_PC_INTERNAL_30 : std_logic ;
  signal CPI_A_INST_INTERNAL : std_logic ;
  signal CPI_A_INST_INTERNAL_0 : std_logic ;
  signal CPI_A_INST_INTERNAL_1 : std_logic ;
  signal CPI_A_INST_INTERNAL_2 : std_logic ;
  signal CPI_A_INST_INTERNAL_3 : std_logic ;
  signal CPI_A_INST_INTERNAL_4 : std_logic ;
  signal CPI_A_INST_INTERNAL_5 : std_logic ;
  signal CPI_A_INST_INTERNAL_6 : std_logic ;
  signal CPI_A_INST_INTERNAL_7 : std_logic ;
  signal CPI_A_INST_INTERNAL_8 : std_logic ;
  signal CPI_A_INST_INTERNAL_9 : std_logic ;
  signal CPI_A_INST_INTERNAL_10 : std_logic ;
  signal CPI_A_INST_INTERNAL_11 : std_logic ;
  signal CPI_A_INST_INTERNAL_12 : std_logic ;
  signal CPI_A_INST_INTERNAL_13 : std_logic ;
  signal CPI_A_INST_INTERNAL_14 : std_logic ;
  signal CPI_A_INST_INTERNAL_15 : std_logic ;
  signal CPI_A_INST_INTERNAL_16 : std_logic ;
  signal CPI_A_INST_INTERNAL_17 : std_logic ;
  signal CPI_A_INST_INTERNAL_18 : std_logic ;
  signal CPI_A_INST_INTERNAL_19 : std_logic ;
  signal CPI_A_INST_INTERNAL_20 : std_logic ;
  signal CPI_A_INST_INTERNAL_21 : std_logic ;
  signal CPI_A_INST_INTERNAL_22 : std_logic ;
  signal CPI_A_INST_INTERNAL_23 : std_logic ;
  signal CPI_A_INST_INTERNAL_24 : std_logic ;
  signal CPI_A_INST_INTERNAL_25 : std_logic ;
  signal CPI_A_INST_INTERNAL_26 : std_logic ;
  signal CPI_A_INST_INTERNAL_27 : std_logic ;
  signal CPI_A_INST_INTERNAL_28 : std_logic ;
  signal CPI_A_INST_INTERNAL_29 : std_logic ;
  signal CPI_A_INST_INTERNAL_30 : std_logic ;
  signal CPI_A_CNT_INTERNAL : std_logic ;
  signal CPI_A_CNT_INTERNAL_0 : std_logic ;
  signal CPI_A_TRAP_INTERNAL : std_logic ;
  signal CPI_A_ANNUL_INTERNAL : std_logic ;
  signal CPI_A_PV_INTERNAL : std_logic ;
  signal CPI_E_PC_INTERNAL : std_logic ;
  signal CPI_E_PC_INTERNAL_0 : std_logic ;
  signal CPI_E_PC_INTERNAL_1 : std_logic ;
  signal CPI_E_PC_INTERNAL_2 : std_logic ;
  signal CPI_E_PC_INTERNAL_3 : std_logic ;
  signal CPI_E_PC_INTERNAL_4 : std_logic ;
  signal CPI_E_PC_INTERNAL_5 : std_logic ;
  signal CPI_E_PC_INTERNAL_6 : std_logic ;
  signal CPI_E_PC_INTERNAL_7 : std_logic ;
  signal CPI_E_PC_INTERNAL_8 : std_logic ;
  signal CPI_E_PC_INTERNAL_9 : std_logic ;
  signal CPI_E_PC_INTERNAL_10 : std_logic ;
  signal CPI_E_PC_INTERNAL_11 : std_logic ;
  signal CPI_E_PC_INTERNAL_12 : std_logic ;
  signal CPI_E_PC_INTERNAL_13 : std_logic ;
  signal CPI_E_PC_INTERNAL_14 : std_logic ;
  signal CPI_E_PC_INTERNAL_15 : std_logic ;
  signal CPI_E_PC_INTERNAL_16 : std_logic ;
  signal CPI_E_PC_INTERNAL_17 : std_logic ;
  signal CPI_E_PC_INTERNAL_18 : std_logic ;
  signal CPI_E_PC_INTERNAL_19 : std_logic ;
  signal CPI_E_PC_INTERNAL_20 : std_logic ;
  signal CPI_E_PC_INTERNAL_21 : std_logic ;
  signal CPI_E_PC_INTERNAL_22 : std_logic ;
  signal CPI_E_PC_INTERNAL_23 : std_logic ;
  signal CPI_E_PC_INTERNAL_24 : std_logic ;
  signal CPI_E_PC_INTERNAL_25 : std_logic ;
  signal CPI_E_PC_INTERNAL_26 : std_logic ;
  signal CPI_E_PC_INTERNAL_27 : std_logic ;
  signal CPI_E_PC_INTERNAL_28 : std_logic ;
  signal CPI_E_PC_INTERNAL_29 : std_logic ;
  signal CPI_E_PC_INTERNAL_30 : std_logic ;
  signal CPI_E_INST_INTERNAL : std_logic ;
  signal CPI_E_INST_INTERNAL_0 : std_logic ;
  signal CPI_E_INST_INTERNAL_1 : std_logic ;
  signal CPI_E_INST_INTERNAL_2 : std_logic ;
  signal CPI_E_INST_INTERNAL_3 : std_logic ;
  signal CPI_E_INST_INTERNAL_4 : std_logic ;
  signal CPI_E_INST_INTERNAL_5 : std_logic ;
  signal CPI_E_INST_INTERNAL_6 : std_logic ;
  signal CPI_E_INST_INTERNAL_7 : std_logic ;
  signal CPI_E_INST_INTERNAL_8 : std_logic ;
  signal CPI_E_INST_INTERNAL_9 : std_logic ;
  signal CPI_E_INST_INTERNAL_10 : std_logic ;
  signal CPI_E_INST_INTERNAL_11 : std_logic ;
  signal CPI_E_INST_INTERNAL_12 : std_logic ;
  signal CPI_E_INST_INTERNAL_13 : std_logic ;
  signal CPI_E_INST_INTERNAL_14 : std_logic ;
  signal CPI_E_INST_INTERNAL_15 : std_logic ;
  signal CPI_E_INST_INTERNAL_16 : std_logic ;
  signal CPI_E_INST_INTERNAL_17 : std_logic ;
  signal CPI_E_INST_INTERNAL_18 : std_logic ;
  signal CPI_E_INST_INTERNAL_19 : std_logic ;
  signal CPI_E_INST_INTERNAL_20 : std_logic ;
  signal CPI_E_INST_INTERNAL_21 : std_logic ;
  signal CPI_E_INST_INTERNAL_22 : std_logic ;
  signal CPI_E_INST_INTERNAL_23 : std_logic ;
  signal CPI_E_INST_INTERNAL_24 : std_logic ;
  signal CPI_E_INST_INTERNAL_25 : std_logic ;
  signal CPI_E_INST_INTERNAL_26 : std_logic ;
  signal CPI_E_INST_INTERNAL_27 : std_logic ;
  signal CPI_E_INST_INTERNAL_28 : std_logic ;
  signal CPI_E_INST_INTERNAL_29 : std_logic ;
  signal CPI_E_INST_INTERNAL_30 : std_logic ;
  signal CPI_E_CNT_INTERNAL : std_logic ;
  signal CPI_E_CNT_INTERNAL_0 : std_logic ;
  signal CPI_E_TRAP_INTERNAL : std_logic ;
  signal CPI_E_ANNUL_INTERNAL : std_logic ;
  signal CPI_E_PV_INTERNAL : std_logic ;
  signal CPI_M_PC_INTERNAL : std_logic ;
  signal CPI_M_PC_INTERNAL_0 : std_logic ;
  signal CPI_M_PC_INTERNAL_1 : std_logic ;
  signal CPI_M_PC_INTERNAL_2 : std_logic ;
  signal CPI_M_PC_INTERNAL_3 : std_logic ;
  signal CPI_M_PC_INTERNAL_4 : std_logic ;
  signal CPI_M_PC_INTERNAL_5 : std_logic ;
  signal CPI_M_PC_INTERNAL_6 : std_logic ;
  signal CPI_M_PC_INTERNAL_7 : std_logic ;
  signal CPI_M_PC_INTERNAL_8 : std_logic ;
  signal CPI_M_PC_INTERNAL_9 : std_logic ;
  signal CPI_M_PC_INTERNAL_10 : std_logic ;
  signal CPI_M_PC_INTERNAL_11 : std_logic ;
  signal CPI_M_PC_INTERNAL_12 : std_logic ;
  signal CPI_M_PC_INTERNAL_13 : std_logic ;
  signal CPI_M_PC_INTERNAL_14 : std_logic ;
  signal CPI_M_PC_INTERNAL_15 : std_logic ;
  signal CPI_M_PC_INTERNAL_16 : std_logic ;
  signal CPI_M_PC_INTERNAL_17 : std_logic ;
  signal CPI_M_PC_INTERNAL_18 : std_logic ;
  signal CPI_M_PC_INTERNAL_19 : std_logic ;
  signal CPI_M_PC_INTERNAL_20 : std_logic ;
  signal CPI_M_PC_INTERNAL_21 : std_logic ;
  signal CPI_M_PC_INTERNAL_22 : std_logic ;
  signal CPI_M_PC_INTERNAL_23 : std_logic ;
  signal CPI_M_PC_INTERNAL_24 : std_logic ;
  signal CPI_M_PC_INTERNAL_25 : std_logic ;
  signal CPI_M_PC_INTERNAL_26 : std_logic ;
  signal CPI_M_PC_INTERNAL_27 : std_logic ;
  signal CPI_M_PC_INTERNAL_28 : std_logic ;
  signal CPI_M_PC_INTERNAL_29 : std_logic ;
  signal CPI_M_PC_INTERNAL_30 : std_logic ;
  signal CPI_M_INST_INTERNAL : std_logic ;
  signal CPI_M_INST_INTERNAL_0 : std_logic ;
  signal CPI_M_INST_INTERNAL_1 : std_logic ;
  signal CPI_M_INST_INTERNAL_2 : std_logic ;
  signal CPI_M_INST_INTERNAL_3 : std_logic ;
  signal CPI_M_INST_INTERNAL_4 : std_logic ;
  signal CPI_M_INST_INTERNAL_5 : std_logic ;
  signal CPI_M_INST_INTERNAL_6 : std_logic ;
  signal CPI_M_INST_INTERNAL_7 : std_logic ;
  signal CPI_M_INST_INTERNAL_8 : std_logic ;
  signal CPI_M_INST_INTERNAL_9 : std_logic ;
  signal CPI_M_INST_INTERNAL_10 : std_logic ;
  signal CPI_M_INST_INTERNAL_11 : std_logic ;
  signal CPI_M_INST_INTERNAL_12 : std_logic ;
  signal CPI_M_INST_INTERNAL_13 : std_logic ;
  signal CPI_M_INST_INTERNAL_14 : std_logic ;
  signal CPI_M_INST_INTERNAL_15 : std_logic ;
  signal CPI_M_INST_INTERNAL_16 : std_logic ;
  signal CPI_M_INST_INTERNAL_17 : std_logic ;
  signal CPI_M_INST_INTERNAL_18 : std_logic ;
  signal CPI_M_INST_INTERNAL_19 : std_logic ;
  signal CPI_M_INST_INTERNAL_20 : std_logic ;
  signal CPI_M_INST_INTERNAL_21 : std_logic ;
  signal CPI_M_INST_INTERNAL_22 : std_logic ;
  signal CPI_M_INST_INTERNAL_23 : std_logic ;
  signal CPI_M_INST_INTERNAL_24 : std_logic ;
  signal CPI_M_INST_INTERNAL_25 : std_logic ;
  signal CPI_M_INST_INTERNAL_26 : std_logic ;
  signal CPI_M_INST_INTERNAL_27 : std_logic ;
  signal CPI_M_INST_INTERNAL_28 : std_logic ;
  signal CPI_M_INST_INTERNAL_29 : std_logic ;
  signal CPI_M_INST_INTERNAL_30 : std_logic ;
  signal CPI_M_CNT_INTERNAL : std_logic ;
  signal CPI_M_CNT_INTERNAL_0 : std_logic ;
  signal CPI_M_TRAP_INTERNAL : std_logic ;
  signal CPI_M_ANNUL_INTERNAL : std_logic ;
  signal CPI_M_PV_INTERNAL : std_logic ;
  signal CPI_X_PC_INTERNAL : std_logic ;
  signal CPI_X_PC_INTERNAL_0 : std_logic ;
  signal CPI_X_PC_INTERNAL_1 : std_logic ;
  signal CPI_X_PC_INTERNAL_2 : std_logic ;
  signal CPI_X_PC_INTERNAL_3 : std_logic ;
  signal CPI_X_PC_INTERNAL_4 : std_logic ;
  signal CPI_X_PC_INTERNAL_5 : std_logic ;
  signal CPI_X_PC_INTERNAL_6 : std_logic ;
  signal CPI_X_PC_INTERNAL_7 : std_logic ;
  signal CPI_X_PC_INTERNAL_8 : std_logic ;
  signal CPI_X_PC_INTERNAL_9 : std_logic ;
  signal CPI_X_PC_INTERNAL_10 : std_logic ;
  signal CPI_X_PC_INTERNAL_11 : std_logic ;
  signal CPI_X_PC_INTERNAL_12 : std_logic ;
  signal CPI_X_PC_INTERNAL_13 : std_logic ;
  signal CPI_X_PC_INTERNAL_14 : std_logic ;
  signal CPI_X_PC_INTERNAL_15 : std_logic ;
  signal CPI_X_PC_INTERNAL_16 : std_logic ;
  signal CPI_X_PC_INTERNAL_17 : std_logic ;
  signal CPI_X_PC_INTERNAL_18 : std_logic ;
  signal CPI_X_PC_INTERNAL_19 : std_logic ;
  signal CPI_X_PC_INTERNAL_20 : std_logic ;
  signal CPI_X_PC_INTERNAL_21 : std_logic ;
  signal CPI_X_PC_INTERNAL_22 : std_logic ;
  signal CPI_X_PC_INTERNAL_23 : std_logic ;
  signal CPI_X_PC_INTERNAL_24 : std_logic ;
  signal CPI_X_PC_INTERNAL_25 : std_logic ;
  signal CPI_X_PC_INTERNAL_26 : std_logic ;
  signal CPI_X_PC_INTERNAL_27 : std_logic ;
  signal CPI_X_PC_INTERNAL_28 : std_logic ;
  signal CPI_X_PC_INTERNAL_29 : std_logic ;
  signal CPI_X_PC_INTERNAL_30 : std_logic ;
  signal CPI_X_INST_INTERNAL : std_logic ;
  signal CPI_X_INST_INTERNAL_0 : std_logic ;
  signal CPI_X_INST_INTERNAL_1 : std_logic ;
  signal CPI_X_INST_INTERNAL_2 : std_logic ;
  signal CPI_X_INST_INTERNAL_3 : std_logic ;
  signal CPI_X_INST_INTERNAL_4 : std_logic ;
  signal CPI_X_INST_INTERNAL_5 : std_logic ;
  signal CPI_X_INST_INTERNAL_6 : std_logic ;
  signal CPI_X_INST_INTERNAL_7 : std_logic ;
  signal CPI_X_INST_INTERNAL_8 : std_logic ;
  signal CPI_X_INST_INTERNAL_9 : std_logic ;
  signal CPI_X_INST_INTERNAL_10 : std_logic ;
  signal CPI_X_INST_INTERNAL_11 : std_logic ;
  signal CPI_X_INST_INTERNAL_12 : std_logic ;
  signal CPI_X_INST_INTERNAL_13 : std_logic ;
  signal CPI_X_INST_INTERNAL_14 : std_logic ;
  signal CPI_X_INST_INTERNAL_15 : std_logic ;
  signal CPI_X_INST_INTERNAL_16 : std_logic ;
  signal CPI_X_INST_INTERNAL_17 : std_logic ;
  signal CPI_X_INST_INTERNAL_18 : std_logic ;
  signal CPI_X_INST_INTERNAL_19 : std_logic ;
  signal CPI_X_INST_INTERNAL_20 : std_logic ;
  signal CPI_X_INST_INTERNAL_21 : std_logic ;
  signal CPI_X_INST_INTERNAL_22 : std_logic ;
  signal CPI_X_INST_INTERNAL_23 : std_logic ;
  signal CPI_X_INST_INTERNAL_24 : std_logic ;
  signal CPI_X_INST_INTERNAL_25 : std_logic ;
  signal CPI_X_INST_INTERNAL_26 : std_logic ;
  signal CPI_X_INST_INTERNAL_27 : std_logic ;
  signal CPI_X_INST_INTERNAL_28 : std_logic ;
  signal CPI_X_INST_INTERNAL_29 : std_logic ;
  signal CPI_X_INST_INTERNAL_30 : std_logic ;
  signal CPI_X_CNT_INTERNAL : std_logic ;
  signal CPI_X_CNT_INTERNAL_0 : std_logic ;
  signal CPI_X_TRAP_INTERNAL : std_logic ;
  signal CPI_X_ANNUL_INTERNAL : std_logic ;
  signal CPI_X_PV_INTERNAL : std_logic ;
  signal CPI_LDDATA_INTERNAL : std_logic ;
  signal CPI_LDDATA_INTERNAL_0 : std_logic ;
  signal CPI_LDDATA_INTERNAL_1 : std_logic ;
  signal CPI_LDDATA_INTERNAL_2 : std_logic ;
  signal CPI_LDDATA_INTERNAL_3 : std_logic ;
  signal CPI_LDDATA_INTERNAL_4 : std_logic ;
  signal CPI_LDDATA_INTERNAL_5 : std_logic ;
  signal CPI_LDDATA_INTERNAL_6 : std_logic ;
  signal CPI_LDDATA_INTERNAL_7 : std_logic ;
  signal CPI_LDDATA_INTERNAL_8 : std_logic ;
  signal CPI_LDDATA_INTERNAL_9 : std_logic ;
  signal CPI_LDDATA_INTERNAL_10 : std_logic ;
  signal CPI_LDDATA_INTERNAL_11 : std_logic ;
  signal CPI_LDDATA_INTERNAL_12 : std_logic ;
  signal CPI_LDDATA_INTERNAL_13 : std_logic ;
  signal CPI_LDDATA_INTERNAL_14 : std_logic ;
  signal CPI_LDDATA_INTERNAL_15 : std_logic ;
  signal CPI_LDDATA_INTERNAL_16 : std_logic ;
  signal CPI_LDDATA_INTERNAL_17 : std_logic ;
  signal CPI_LDDATA_INTERNAL_18 : std_logic ;
  signal CPI_LDDATA_INTERNAL_19 : std_logic ;
  signal CPI_LDDATA_INTERNAL_20 : std_logic ;
  signal CPI_LDDATA_INTERNAL_21 : std_logic ;
  signal CPI_LDDATA_INTERNAL_22 : std_logic ;
  signal CPI_LDDATA_INTERNAL_23 : std_logic ;
  signal CPI_LDDATA_INTERNAL_24 : std_logic ;
  signal CPI_LDDATA_INTERNAL_25 : std_logic ;
  signal CPI_LDDATA_INTERNAL_26 : std_logic ;
  signal CPI_LDDATA_INTERNAL_27 : std_logic ;
  signal CPI_LDDATA_INTERNAL_28 : std_logic ;
  signal CPI_LDDATA_INTERNAL_29 : std_logic ;
  signal CPI_LDDATA_INTERNAL_30 : std_logic ;
  signal CPI_DBG_ENABLE_INTERNAL : std_logic ;
  signal CPI_DBG_WRITE_INTERNAL : std_logic ;
  signal CPI_DBG_FSR_INTERNAL : std_logic ;
  signal CPI_DBG_ADDR_INTERNAL : std_logic ;
  signal CPI_DBG_ADDR_INTERNAL_0 : std_logic ;
  signal CPI_DBG_ADDR_INTERNAL_1 : std_logic ;
  signal CPI_DBG_ADDR_INTERNAL_2 : std_logic ;
  signal CPI_DBG_ADDR_INTERNAL_3 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_0 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_1 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_2 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_3 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_4 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_5 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_6 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_7 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_8 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_9 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_10 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_11 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_12 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_13 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_14 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_15 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_16 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_17 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_18 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_19 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_20 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_21 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_22 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_23 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_24 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_25 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_26 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_27 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_28 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_29 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_30 : std_logic ;
  signal RFO1_DATA1_INTERNAL : std_logic ;
  signal RFO1_DATA1_INTERNAL_0 : std_logic ;
  signal RFO1_DATA1_INTERNAL_1 : std_logic ;
  signal RFO1_DATA1_INTERNAL_2 : std_logic ;
  signal RFO1_DATA1_INTERNAL_3 : std_logic ;
  signal RFO1_DATA1_INTERNAL_4 : std_logic ;
  signal RFO1_DATA1_INTERNAL_5 : std_logic ;
  signal RFO1_DATA1_INTERNAL_6 : std_logic ;
  signal RFO1_DATA1_INTERNAL_7 : std_logic ;
  signal RFO1_DATA1_INTERNAL_8 : std_logic ;
  signal RFO1_DATA1_INTERNAL_9 : std_logic ;
  signal RFO1_DATA1_INTERNAL_10 : std_logic ;
  signal RFO1_DATA1_INTERNAL_11 : std_logic ;
  signal RFO1_DATA1_INTERNAL_12 : std_logic ;
  signal RFO1_DATA1_INTERNAL_13 : std_logic ;
  signal RFO1_DATA1_INTERNAL_14 : std_logic ;
  signal RFO1_DATA1_INTERNAL_15 : std_logic ;
  signal RFO1_DATA1_INTERNAL_16 : std_logic ;
  signal RFO1_DATA1_INTERNAL_17 : std_logic ;
  signal RFO1_DATA1_INTERNAL_18 : std_logic ;
  signal RFO1_DATA1_INTERNAL_19 : std_logic ;
  signal RFO1_DATA1_INTERNAL_20 : std_logic ;
  signal RFO1_DATA1_INTERNAL_21 : std_logic ;
  signal RFO1_DATA1_INTERNAL_22 : std_logic ;
  signal RFO1_DATA1_INTERNAL_23 : std_logic ;
  signal RFO1_DATA1_INTERNAL_24 : std_logic ;
  signal RFO1_DATA1_INTERNAL_25 : std_logic ;
  signal RFO1_DATA1_INTERNAL_26 : std_logic ;
  signal RFO1_DATA1_INTERNAL_27 : std_logic ;
  signal RFO1_DATA1_INTERNAL_28 : std_logic ;
  signal RFO1_DATA1_INTERNAL_29 : std_logic ;
  signal RFO1_DATA1_INTERNAL_30 : std_logic ;
  signal RFO1_DATA2_INTERNAL : std_logic ;
  signal RFO1_DATA2_INTERNAL_0 : std_logic ;
  signal RFO1_DATA2_INTERNAL_1 : std_logic ;
  signal RFO1_DATA2_INTERNAL_2 : std_logic ;
  signal RFO1_DATA2_INTERNAL_3 : std_logic ;
  signal RFO1_DATA2_INTERNAL_4 : std_logic ;
  signal RFO1_DATA2_INTERNAL_5 : std_logic ;
  signal RFO1_DATA2_INTERNAL_6 : std_logic ;
  signal RFO1_DATA2_INTERNAL_7 : std_logic ;
  signal RFO1_DATA2_INTERNAL_8 : std_logic ;
  signal RFO1_DATA2_INTERNAL_9 : std_logic ;
  signal RFO1_DATA2_INTERNAL_10 : std_logic ;
  signal RFO1_DATA2_INTERNAL_11 : std_logic ;
  signal RFO1_DATA2_INTERNAL_12 : std_logic ;
  signal RFO1_DATA2_INTERNAL_13 : std_logic ;
  signal RFO1_DATA2_INTERNAL_14 : std_logic ;
  signal RFO1_DATA2_INTERNAL_15 : std_logic ;
  signal RFO1_DATA2_INTERNAL_16 : std_logic ;
  signal RFO1_DATA2_INTERNAL_17 : std_logic ;
  signal RFO1_DATA2_INTERNAL_18 : std_logic ;
  signal RFO1_DATA2_INTERNAL_19 : std_logic ;
  signal RFO1_DATA2_INTERNAL_20 : std_logic ;
  signal RFO1_DATA2_INTERNAL_21 : std_logic ;
  signal RFO1_DATA2_INTERNAL_22 : std_logic ;
  signal RFO1_DATA2_INTERNAL_23 : std_logic ;
  signal RFO1_DATA2_INTERNAL_24 : std_logic ;
  signal RFO1_DATA2_INTERNAL_25 : std_logic ;
  signal RFO1_DATA2_INTERNAL_26 : std_logic ;
  signal RFO1_DATA2_INTERNAL_27 : std_logic ;
  signal RFO1_DATA2_INTERNAL_28 : std_logic ;
  signal RFO1_DATA2_INTERNAL_29 : std_logic ;
  signal RFO1_DATA2_INTERNAL_30 : std_logic ;
  signal RFO2_DATA1_INTERNAL : std_logic ;
  signal RFO2_DATA1_INTERNAL_0 : std_logic ;
  signal RFO2_DATA1_INTERNAL_1 : std_logic ;
  signal RFO2_DATA1_INTERNAL_2 : std_logic ;
  signal RFO2_DATA1_INTERNAL_3 : std_logic ;
  signal RFO2_DATA1_INTERNAL_4 : std_logic ;
  signal RFO2_DATA1_INTERNAL_5 : std_logic ;
  signal RFO2_DATA1_INTERNAL_6 : std_logic ;
  signal RFO2_DATA1_INTERNAL_7 : std_logic ;
  signal RFO2_DATA1_INTERNAL_8 : std_logic ;
  signal RFO2_DATA1_INTERNAL_9 : std_logic ;
  signal RFO2_DATA1_INTERNAL_10 : std_logic ;
  signal RFO2_DATA1_INTERNAL_11 : std_logic ;
  signal RFO2_DATA1_INTERNAL_12 : std_logic ;
  signal RFO2_DATA1_INTERNAL_13 : std_logic ;
  signal RFO2_DATA1_INTERNAL_14 : std_logic ;
  signal RFO2_DATA1_INTERNAL_15 : std_logic ;
  signal RFO2_DATA1_INTERNAL_16 : std_logic ;
  signal RFO2_DATA1_INTERNAL_17 : std_logic ;
  signal RFO2_DATA1_INTERNAL_18 : std_logic ;
  signal RFO2_DATA1_INTERNAL_19 : std_logic ;
  signal RFO2_DATA1_INTERNAL_20 : std_logic ;
  signal RFO2_DATA1_INTERNAL_21 : std_logic ;
  signal RFO2_DATA1_INTERNAL_22 : std_logic ;
  signal RFO2_DATA1_INTERNAL_23 : std_logic ;
  signal RFO2_DATA1_INTERNAL_24 : std_logic ;
  signal RFO2_DATA1_INTERNAL_25 : std_logic ;
  signal RFO2_DATA1_INTERNAL_26 : std_logic ;
  signal RFO2_DATA1_INTERNAL_27 : std_logic ;
  signal RFO2_DATA1_INTERNAL_28 : std_logic ;
  signal RFO2_DATA1_INTERNAL_29 : std_logic ;
  signal RFO2_DATA1_INTERNAL_30 : std_logic ;
  signal RFO2_DATA2_INTERNAL : std_logic ;
  signal RFO2_DATA2_INTERNAL_0 : std_logic ;
  signal RFO2_DATA2_INTERNAL_1 : std_logic ;
  signal RFO2_DATA2_INTERNAL_2 : std_logic ;
  signal RFO2_DATA2_INTERNAL_3 : std_logic ;
  signal RFO2_DATA2_INTERNAL_4 : std_logic ;
  signal RFO2_DATA2_INTERNAL_5 : std_logic ;
  signal RFO2_DATA2_INTERNAL_6 : std_logic ;
  signal RFO2_DATA2_INTERNAL_7 : std_logic ;
  signal RFO2_DATA2_INTERNAL_8 : std_logic ;
  signal RFO2_DATA2_INTERNAL_9 : std_logic ;
  signal RFO2_DATA2_INTERNAL_10 : std_logic ;
  signal RFO2_DATA2_INTERNAL_11 : std_logic ;
  signal RFO2_DATA2_INTERNAL_12 : std_logic ;
  signal RFO2_DATA2_INTERNAL_13 : std_logic ;
  signal RFO2_DATA2_INTERNAL_14 : std_logic ;
  signal RFO2_DATA2_INTERNAL_15 : std_logic ;
  signal RFO2_DATA2_INTERNAL_16 : std_logic ;
  signal RFO2_DATA2_INTERNAL_17 : std_logic ;
  signal RFO2_DATA2_INTERNAL_18 : std_logic ;
  signal RFO2_DATA2_INTERNAL_19 : std_logic ;
  signal RFO2_DATA2_INTERNAL_20 : std_logic ;
  signal RFO2_DATA2_INTERNAL_21 : std_logic ;
  signal RFO2_DATA2_INTERNAL_22 : std_logic ;
  signal RFO2_DATA2_INTERNAL_23 : std_logic ;
  signal RFO2_DATA2_INTERNAL_24 : std_logic ;
  signal RFO2_DATA2_INTERNAL_25 : std_logic ;
  signal RFO2_DATA2_INTERNAL_26 : std_logic ;
  signal RFO2_DATA2_INTERNAL_27 : std_logic ;
  signal RFO2_DATA2_INTERNAL_28 : std_logic ;
  signal RFO2_DATA2_INTERNAL_29 : std_logic ;
  signal RFO2_DATA2_INTERNAL_30 : std_logic ;
  signal VCC : std_logic ;
  signal GND : std_logic ;
  signal \GRLFPC2_0.FPI.START\ : std_logic ;
  signal \GRLFPC2_0.FPI.RST\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\ : std_logic ;
  signal \GRLFPC2_0.R.I.EXEC\ : std_logic ;
  signal \GRLFPC2_0.R.X.LD\ : std_logic ;
  signal \GRLFPC2_0.R.X.AFSR\ : std_logic ;
  signal \GRLFPC2_0.R.X.SEQERR\ : std_logic ;
  signal \GRLFPC2_0.R.X.FPOP\ : std_logic ;
  signal \GRLFPC2_0.R.MK.HOLDN1\ : std_logic ;
  signal \GRLFPC2_0.R.E.FPOP\ : std_logic ;
  signal \GRLFPC2_0.R.M.FPOP\ : std_logic ;
  signal \GRLFPC2_0.R.MK.HOLDN2\ : std_logic ;
  signal \GRLFPC2_0.R.I.V\ : std_logic ;
  signal \GRLFPC2_0.R.M.LD\ : std_logic ;
  signal \GRLFPC2_0.R.E.LD\ : std_logic ;
  signal \GRLFPC2_0.R.A.LD\ : std_logic ;
  signal \GRLFPC2_0.R.A.FPOP\ : std_logic ;
  signal \GRLFPC2_0.R.X.AFQ\ : std_logic ;
  signal \GRLFPC2_0.R.I.RDD\ : std_logic ;
  signal \GRLFPC2_0.R.X.RDD\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.NONSTD\ : std_logic ;
  signal \GRLFPC2_0.N_554\ : std_logic ;
  signal \GRLFPC2_0.N_557\ : std_logic ;
  signal \GRLFPC2_0.N_558\ : std_logic ;
  signal \GRLFPC2_0.N_559\ : std_logic ;
  signal \GRLFPC2_0.R.MK.RST2\ : std_logic ;
  signal \GRLFPC2_0.R.MK.RST\ : std_logic ;
  signal \GRLFPC2_0.R.A.RS1D\ : std_logic ;
  signal \GRLFPC2_0.R.A.RS2D\ : std_logic ;
  signal \GRLFPC2_0.N_553\ : std_logic ;
  signal \GRLFPC2_0.R.E.AFQ_O\ : std_logic ;
  signal \GRLFPC2_0.N_1829_O\ : std_logic ;
  signal \GRLFPC2_0.R.E.AFSR_O\ : std_logic ;
  signal \GRLFPC2_0.R.A.AFQ_O\ : std_logic ;
  signal \GRLFPC2_0.R.A.AFSR_O\ : std_logic ;
  signal \GRLFPC2_0.COMB.LOCKGEN.LOCKI_O\ : std_logic ;
  signal \GRLFPC2_0.COMB.FPDECODE.ST_O\ : std_logic ;
  signal \GRLFPC2_0.HOLDN_O\ : std_logic ;
  signal \GRLFPC2_0.COMB.LOCKGEN.LOCKI_O_3\ : std_logic ;
  signal \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\ : std_logic ;
  signal \GRLFPC2_0.COMB.ANNULFPU_1_O\ : std_logic ;
  signal \GRLFPC2_0.R.MK.RST2_O\ : std_logic ;
  signal \GRLFPC2_0.R.MK.HOLDN2_O\ : std_logic ;
  signal \GRLFPC2_0.R.MK.HOLDN1_O_0\ : std_logic ;
  signal \GRLFPC2_0.R.MK.HOLDN2_O_0\ : std_logic ;
  signal \GRLFPC2_0.R.MK.RST_O_0\ : std_logic ;
  signal \GRLFPC2_0.R.MK.RST2_O_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.ANNULFPU_1_O_0\ : std_logic ;
  signal \GRLFPC2_0.R.MK.BUSY_O\ : std_logic ;
  signal \GRLFPC2_0.N_1837_O\ : std_logic ;
  signal \GRLFPC2_0.N_95\ : std_logic ;
  signal \GRLFPC2_0.N_96\ : std_logic ;
  signal \GRLFPC2_0.N_97\ : std_logic ;
  signal \GRLFPC2_0.N_98\ : std_logic ;
  signal \GRLFPC2_0.N_99\ : std_logic ;
  signal \GRLFPC2_0.N_100\ : std_logic ;
  signal \GRLFPC2_0.N_101\ : std_logic ;
  signal \GRLFPC2_0.N_102\ : std_logic ;
  signal \GRLFPC2_0.N_103\ : std_logic ;
  signal \GRLFPC2_0.N_104\ : std_logic ;
  signal \GRLFPC2_0.N_105\ : std_logic ;
  signal \GRLFPC2_0.N_106\ : std_logic ;
  signal \GRLFPC2_0.N_107\ : std_logic ;
  signal \GRLFPC2_0.N_108\ : std_logic ;
  signal \GRLFPC2_0.N_109\ : std_logic ;
  signal \GRLFPC2_0.N_110\ : std_logic ;
  signal \GRLFPC2_0.N_111\ : std_logic ;
  signal \GRLFPC2_0.N_112\ : std_logic ;
  signal \GRLFPC2_0.N_113\ : std_logic ;
  signal \GRLFPC2_0.N_114\ : std_logic ;
  signal \GRLFPC2_0.N_115\ : std_logic ;
  signal \GRLFPC2_0.N_116\ : std_logic ;
  signal \GRLFPC2_0.N_117\ : std_logic ;
  signal \GRLFPC2_0.N_118\ : std_logic ;
  signal \GRLFPC2_0.N_119\ : std_logic ;
  signal \GRLFPC2_0.N_120\ : std_logic ;
  signal \GRLFPC2_0.N_121\ : std_logic ;
  signal \GRLFPC2_0.N_122\ : std_logic ;
  signal \GRLFPC2_0.N_123\ : std_logic ;
  signal \GRLFPC2_0.N_124\ : std_logic ;
  signal \GRLFPC2_0.N_125\ : std_logic ;
  signal \GRLFPC2_0.N_126\ : std_logic ;
  signal \GRLFPC2_0.N_127\ : std_logic ;
  signal \GRLFPC2_0.N_128\ : std_logic ;
  signal \GRLFPC2_0.N_129\ : std_logic ;
  signal \GRLFPC2_0.N_130\ : std_logic ;
  signal \GRLFPC2_0.N_131\ : std_logic ;
  signal \GRLFPC2_0.N_132\ : std_logic ;
  signal \GRLFPC2_0.N_133\ : std_logic ;
  signal \GRLFPC2_0.N_134\ : std_logic ;
  signal \GRLFPC2_0.N_135\ : std_logic ;
  signal \GRLFPC2_0.N_136\ : std_logic ;
  signal \GRLFPC2_0.N_137\ : std_logic ;
  signal \GRLFPC2_0.N_2103\ : std_logic ;
  signal \GRLFPC2_0.N_2105\ : std_logic ;
  signal \GRLFPC2_0.N_2111\ : std_logic ;
  signal \GRLFPC2_0.COMB.ANNULFPU_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.RS1D_1\ : std_logic ;
  signal \GRLFPC2_0.N_3150\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5410\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5391\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN25_NOTPROP\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_954\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4459\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4874\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7259\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7260\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7272\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7274\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10017\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10018\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10019\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10020\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10021\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10022\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10023\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10024\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10025\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10026\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10027\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10028\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10029\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10030\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10031\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10032\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10033\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10034\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10035\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10036\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10037\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10038\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10039\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10040\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10041\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10042\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10043\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10044\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10045\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10046\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10047\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10048\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10049\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10050\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10051\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10052\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10053\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10054\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10055\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10056\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10061\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10064\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10066\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10067\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10069\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10070\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10071\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10072\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10074\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10077\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10078\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10079\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10080\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10081\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10082\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10084\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10085\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10086\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10087\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10088\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10089\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10090\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10091\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10092\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10093\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10094\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10095\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10096\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10097\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10098\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10099\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10100\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10101\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10102\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10103\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10104\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10105\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10106\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10107\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10108\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10109\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10110\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10111\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10112\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10113\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10114\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10115\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10116\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10117\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10118\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10119\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10120\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10121\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10122\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10123\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10124\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10125\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10126\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10127\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10128\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10129\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10130\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10131\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10132\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10133\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10134\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10552\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SFTLFT.AREGXORBREG\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3926\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_770\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_551\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_479\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1809\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1758\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_513\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1769\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_812\ : std_logic ;
  signal N_1 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.UN36_PCTRL_NEW_I\ : std_logic ;
  signal N_27258 : std_logic ;
  signal N_27259 : std_logic ;
  signal N_27260 : std_logic ;
  signal N_27261 : std_logic ;
  signal N_27262 : std_logic ;
  signal N_27263 : std_logic ;
  signal N_27264 : std_logic ;
  signal N_27265 : std_logic ;
  signal N_27266 : std_logic ;
  signal N_27267 : std_logic ;
  signal N_27268 : std_logic ;
  signal N_27269 : std_logic ;
  signal N_27270 : std_logic ;
  signal N_27271 : std_logic ;
  signal N_27272 : std_logic ;
  signal N_27273 : std_logic ;
  signal N_27274 : std_logic ;
  signal N_27275 : std_logic ;
  signal N_27276 : std_logic ;
  signal N_27277 : std_logic ;
  signal N_27278 : std_logic ;
  signal N_27279 : std_logic ;
  signal N_27280 : std_logic ;
  signal N_27281 : std_logic ;
  signal N_27282 : std_logic ;
  signal N_27283 : std_logic ;
  signal N_27284 : std_logic ;
  signal N_27285 : std_logic ;
  signal N_27286 : std_logic ;
  signal N_27287 : std_logic ;
  signal N_27288 : std_logic ;
  signal N_27289 : std_logic ;
  signal N_27290 : std_logic ;
  signal N_27291 : std_logic ;
  signal N_27292 : std_logic ;
  signal N_27293 : std_logic ;
  signal N_27294 : std_logic ;
  signal N_27295 : std_logic ;
  signal N_27296 : std_logic ;
  signal N_27297 : std_logic ;
  signal N_27298 : std_logic ;
  signal N_27299 : std_logic ;
  signal N_27300 : std_logic ;
  signal N_27301 : std_logic ;
  signal N_27302 : std_logic ;
  signal N_27303 : std_logic ;
  signal N_27304 : std_logic ;
  signal N_27305 : std_logic ;
  signal N_27306 : std_logic ;
  signal N_27307 : std_logic ;
  signal N_27308 : std_logic ;
  signal N_27309 : std_logic ;
  signal N_27310 : std_logic ;
  signal N_27311 : std_logic ;
  signal N_27312 : std_logic ;
  signal N_27313 : std_logic ;
  signal N_27314 : std_logic ;
  signal N_27315 : std_logic ;
  signal N_27316 : std_logic ;
  signal N_29683 : std_logic ;
  signal N_29684 : std_logic ;
  signal N_29686 : std_logic ;
  signal N_29687 : std_logic ;
  signal N_29689 : std_logic ;
  signal N_29690 : std_logic ;
  signal N_29692 : std_logic ;
  signal N_29693 : std_logic ;
  signal N_29695 : std_logic ;
  signal N_29696 : std_logic ;
  signal N_29698 : std_logic ;
  signal N_29699 : std_logic ;
  signal N_29701 : std_logic ;
  signal N_29702 : std_logic ;
  signal N_29704 : std_logic ;
  signal N_29705 : std_logic ;
  signal N_29707 : std_logic ;
  signal N_29708 : std_logic ;
  signal N_29710 : std_logic ;
  signal N_29711 : std_logic ;
  signal N_29713 : std_logic ;
  signal N_29714 : std_logic ;
  signal N_29716 : std_logic ;
  signal N_29717 : std_logic ;
  signal N_29719 : std_logic ;
  signal N_29720 : std_logic ;
  signal N_29722 : std_logic ;
  signal N_29723 : std_logic ;
  signal N_29725 : std_logic ;
  signal N_29726 : std_logic ;
  signal N_29728 : std_logic ;
  signal N_29729 : std_logic ;
  signal N_29731 : std_logic ;
  signal N_29732 : std_logic ;
  signal N_29734 : std_logic ;
  signal N_29735 : std_logic ;
  signal N_29737 : std_logic ;
  signal N_29738 : std_logic ;
  signal N_29740 : std_logic ;
  signal N_29741 : std_logic ;
  signal N_29743 : std_logic ;
  signal N_29744 : std_logic ;
  signal N_29746 : std_logic ;
  signal N_29747 : std_logic ;
  signal N_29749 : std_logic ;
  signal N_29750 : std_logic ;
  signal N_29752 : std_logic ;
  signal N_29753 : std_logic ;
  signal N_29755 : std_logic ;
  signal N_29756 : std_logic ;
  signal N_29758 : std_logic ;
  signal N_29759 : std_logic ;
  signal N_29761 : std_logic ;
  signal N_29762 : std_logic ;
  signal N_29764 : std_logic ;
  signal N_29765 : std_logic ;
  signal N_29767 : std_logic ;
  signal N_29768 : std_logic ;
  signal N_29770 : std_logic ;
  signal N_29771 : std_logic ;
  signal N_29773 : std_logic ;
  signal N_29774 : std_logic ;
  signal N_29776 : std_logic ;
  signal N_29777 : std_logic ;
  signal N_29779 : std_logic ;
  signal N_29780 : std_logic ;
  signal N_29782 : std_logic ;
  signal N_29783 : std_logic ;
  signal N_29785 : std_logic ;
  signal N_29786 : std_logic ;
  signal N_29788 : std_logic ;
  signal N_29789 : std_logic ;
  signal N_29791 : std_logic ;
  signal N_29792 : std_logic ;
  signal N_29794 : std_logic ;
  signal N_29795 : std_logic ;
  signal N_29797 : std_logic ;
  signal N_29798 : std_logic ;
  signal N_29800 : std_logic ;
  signal N_29801 : std_logic ;
  signal N_29803 : std_logic ;
  signal N_29804 : std_logic ;
  signal N_29806 : std_logic ;
  signal N_29807 : std_logic ;
  signal N_29809 : std_logic ;
  signal N_29810 : std_logic ;
  signal N_29812 : std_logic ;
  signal N_29813 : std_logic ;
  signal N_29815 : std_logic ;
  signal N_29816 : std_logic ;
  signal N_29818 : std_logic ;
  signal N_29819 : std_logic ;
  signal N_29821 : std_logic ;
  signal N_29822 : std_logic ;
  signal N_29824 : std_logic ;
  signal N_29825 : std_logic ;
  signal N_29827 : std_logic ;
  signal N_29828 : std_logic ;
  signal N_29830 : std_logic ;
  signal N_29831 : std_logic ;
  signal N_29833 : std_logic ;
  signal N_29834 : std_logic ;
  signal N_29836 : std_logic ;
  signal N_29837 : std_logic ;
  signal N_29839 : std_logic ;
  signal N_29840 : std_logic ;
  signal N_29842 : std_logic ;
  signal N_29843 : std_logic ;
  signal N_29845 : std_logic ;
  signal N_29846 : std_logic ;
  signal N_29848 : std_logic ;
  signal N_29849 : std_logic ;
  signal N_29851 : std_logic ;
  signal N_29852 : std_logic ;
  signal N_29854 : std_logic ;
  signal N_29855 : std_logic ;
  signal N_29857 : std_logic ;
  signal N_29858 : std_logic ;
  signal N_29860 : std_logic ;
  signal N_29861 : std_logic ;
  signal N_29863 : std_logic ;
  signal N_29864 : std_logic ;
  signal N_29866 : std_logic ;
  signal N_29867 : std_logic ;
  signal N_29869 : std_logic ;
  signal N_29870 : std_logic ;
  signal N_29872 : std_logic ;
  signal N_29873 : std_logic ;
  signal N_29875 : std_logic ;
  signal N_29876 : std_logic ;
  signal N_29878 : std_logic ;
  signal N_29879 : std_logic ;
  signal N_29881 : std_logic ;
  signal N_29882 : std_logic ;
  signal N_29884 : std_logic ;
  signal N_29885 : std_logic ;
  signal N_29887 : std_logic ;
  signal N_29888 : std_logic ;
  signal N_29890 : std_logic ;
  signal N_29891 : std_logic ;
  signal N_29893 : std_logic ;
  signal N_29894 : std_logic ;
  signal N_29896 : std_logic ;
  signal N_29897 : std_logic ;
  signal N_29899 : std_logic ;
  signal N_29900 : std_logic ;
  signal N_29902 : std_logic ;
  signal N_29903 : std_logic ;
  signal N_29905 : std_logic ;
  signal N_29906 : std_logic ;
  signal N_29908 : std_logic ;
  signal N_29909 : std_logic ;
  signal N_29911 : std_logic ;
  signal N_29912 : std_logic ;
  signal N_29914 : std_logic ;
  signal N_29915 : std_logic ;
  signal N_29917 : std_logic ;
  signal N_29918 : std_logic ;
  signal N_29920 : std_logic ;
  signal N_29921 : std_logic ;
  signal N_29923 : std_logic ;
  signal N_29924 : std_logic ;
  signal N_29926 : std_logic ;
  signal N_29927 : std_logic ;
  signal N_29929 : std_logic ;
  signal N_29930 : std_logic ;
  signal N_29932 : std_logic ;
  signal N_29933 : std_logic ;
  signal N_29935 : std_logic ;
  signal N_29936 : std_logic ;
  signal N_29938 : std_logic ;
  signal N_29939 : std_logic ;
  signal N_29941 : std_logic ;
  signal N_29942 : std_logic ;
  signal N_29944 : std_logic ;
  signal N_29945 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6.Z_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6.Z_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6.Z_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_47__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_46__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_44__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_41__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_40__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_39__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_35__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_30__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_24__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_23__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_22__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_21__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_20__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_16__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_15__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_14__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_8__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_2__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_1__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_372__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_319__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_318__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_317__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_316__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_258__N_5_I\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_176__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_175__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_17__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_16__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_15__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_14__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_13__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_12__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_11__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_10__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_9__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_8__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_7__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_6__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_5__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_4__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_3__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_2__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_1__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_0__G2\ : std_logic ;
  signal \GRLFPC2_0.COMB.FPDECODE.ST\ : std_logic ;
  signal \GRLFPC2_0.R.M.AFSR_RET_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.M.AFQ_RET_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.SEQERR_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.COMB.RS2D_1\ : std_logic ;
  signal \GRLFPC2_0.R.A.RDD_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.A.LD_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.A.FPOP_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.FTT_0_0_2__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.FTT_0_0_0__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.NONSTD_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.X.LD_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.X.FPOP_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.X.AFSR_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.X.AFQ_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.M.LD_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.M.FPOP_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.LD_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.E.FPOP_1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_0__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_1__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_2__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_3__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_4__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_5__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_6__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_7__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_8__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_9__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_10__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_11__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_12__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_13__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_14__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_15__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_16__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_17__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_18__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_19__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_20__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_21__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_22__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_23__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_24__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_25__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_26__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_27__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_28__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_29__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_30__G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.STDATA_1_0_31__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.RD_0_0_0__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.RD_0_0_1__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.TEM_1_0_0__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.TEM_1_0_1__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.TEM_1_0_2__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.TEM_1_0_3__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.TEM_1_0_4__G1\ : std_logic ;
  signal \GRLFPC2_0.R.STATE_0_0_0__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.FCC_0_0_0__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.FCC_0_0_1__G1\ : std_logic ;
  signal \GRLFPC2_0.R.I.CC_0_0_0__G2\ : std_logic ;
  signal \GRLFPC2_0.R.I.CC_0_0_1__G2\ : std_logic ;
  signal \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\ : std_logic ;
  signal \GRLFPC2_0.R.I.EXC_2_0_1__G2\ : std_logic ;
  signal \GRLFPC2_0.R.I.EXC_2_0_2__G2\ : std_logic ;
  signal \GRLFPC2_0.R.I.EXC_2_0_3__G2\ : std_logic ;
  signal \GRLFPC2_0.R.I.EXC_2_0_4__G2\ : std_logic ;
  signal N_36985 : std_logic ;
  signal N_36986 : std_logic ;
  signal N_37176 : std_logic ;
  signal N_37203 : std_logic ;
  signal N_37230 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_49_I\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_51_I\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__I0_I_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_48__I0_I_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_11__I0_I_1\ : std_logic ;
  signal N_37415 : std_logic ;
  signal N_37416 : std_logic ;
  signal N_37417 : std_logic ;
  signal N_37418 : std_logic ;
  signal N_37419 : std_logic ;
  signal N_37420 : std_logic ;
  signal N_37421 : std_logic ;
  signal N_37422 : std_logic ;
  signal N_37423 : std_logic ;
  signal N_37424 : std_logic ;
  signal \GRLFPC2_0.N_76_I\ : std_logic ;
  signal N_37428 : std_logic ;
  signal N_37429 : std_logic ;
  signal \GRLFPC2_0.R.STATE_0_0_1__I0_I_1\ : std_logic ;
  signal N_37431 : std_logic ;
  signal N_37432 : std_logic ;
  signal N_37433 : std_logic ;
  signal \GRLFPC2_0.R.FSR.AEXC_1_0_0__I0_I_0\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.AEXC_1_0_1__I0_I_1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.AEXC_1_0_2__I0_I_0\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.AEXC_1_0_3__I0_I_1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.AEXC_1_0_4__I0_I_0\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.CEXC_1_0_0__I0_I_1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.CEXC_1_0_1__I0_I_0\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.CEXC_1_0_2__I0_I_1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.CEXC_1_0_3__I0_I_0\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.CEXC_1_0_4__I0_I_1\ : std_logic ;
  signal N_38487 : std_logic ;
  signal N_38488 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_877_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10911\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10905\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9598\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1736\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11641\ : std_logic ;
  signal N_32831 : std_logic ;
  signal N_34255 : std_logic ;
  signal N_32848 : std_logic ;
  signal N_32838 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_809\ : std_logic ;
  signal N_32821 : std_logic ;
  signal N_28857_1 : std_logic ;
  signal N_33004 : std_logic ;
  signal N_33146_1 : std_logic ;
  signal N_28492_1 : std_logic ;
  signal N_34341_1 : std_logic ;
  signal N_32858_1 : std_logic ;
  signal N_32859_1 : std_logic ;
  signal N_28212_1 : std_logic ;
  signal N_32818_I : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_604\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_603\ : std_logic ;
  signal N_33984_2 : std_logic ;
  signal N_28549_1 : std_logic ;
  signal N_33111 : std_logic ;
  signal N_33179 : std_logic ;
  signal N_33193 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_782\ : std_logic ;
  signal N_33899 : std_logic ;
  signal N_33904 : std_logic ;
  signal N_33134 : std_logic ;
  signal N_33130 : std_logic ;
  signal N_33139 : std_logic ;
  signal N_32978 : std_logic ;
  signal N_32722_2 : std_logic ;
  signal N_32722_1 : std_logic ;
  signal N_29071_1 : std_logic ;
  signal N_28634_1 : std_logic ;
  signal N_32979_1 : std_logic ;
  signal N_33297_1 : std_logic ;
  signal N_32909_1 : std_logic ;
  signal N_33175 : std_logic ;
  signal N_33138_1 : std_logic ;
  signal N_28271_1 : std_logic ;
  signal N_33152_2 : std_logic ;
  signal N_32730_1 : std_logic ;
  signal N_33903 : std_logic ;
  signal N_29195_1 : std_logic ;
  signal N_33574_1 : std_logic ;
  signal N_33607_1 : std_logic ;
  signal N_33543 : std_logic ;
  signal N_29366_1 : std_logic ;
  signal N_28250_1 : std_logic ;
  signal N_29653_1 : std_logic ;
  signal N_29262_1 : std_logic ;
  signal N_34051 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1730\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_458\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_426\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1566\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_475\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9509\ : std_logic ;
  signal N_28266_2 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9514\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1607\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9566\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1757\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_648\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_814\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_816\ : std_logic ;
  signal N_33010 : std_logic ;
  signal N_34056 : std_logic ;
  signal N_34052 : std_logic ;
  signal N_34049 : std_logic ;
  signal N_32723_1 : std_logic ;
  signal N_34055_2 : std_logic ;
  signal N_28564_2 : std_logic ;
  signal N_32782_1 : std_logic ;
  signal N_32738_2 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5330\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8524\ : std_logic ;
  signal N_28264_1 : std_logic ;
  signal N_29518_1 : std_logic ;
  signal N_32982_1 : std_logic ;
  signal N_33276 : std_logic ;
  signal N_28261_1 : std_logic ;
  signal N_28222_1 : std_logic ;
  signal N_33548 : std_logic ;
  signal N_33178 : std_logic ;
  signal N_33411 : std_logic ;
  signal N_34233 : std_logic ;
  signal N_33436_1 : std_logic ;
  signal N_32796_2 : std_logic ;
  signal N_33023 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9418\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_544\ : std_logic ;
  signal N_33445 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1304\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9158\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8764\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_769\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9200\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9159\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_659\ : std_logic ;
  signal N_34334 : std_logic ;
  signal N_33499 : std_logic ;
  signal N_32899 : std_logic ;
  signal N_33207 : std_logic ;
  signal N_33916 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1055\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9165\ : std_logic ;
  signal N_33081_1 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1659\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9502\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1237\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9503\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_797\ : std_logic ;
  signal N_33577_1 : std_logic ;
  signal N_28243 : std_logic ;
  signal N_33659_1 : std_logic ;
  signal N_28560_2 : std_logic ;
  signal N_28210 : std_logic ;
  signal N_32844_3 : std_logic ;
  signal N_28208_2 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9369\ : std_logic ;
  signal N_33798_I : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1187\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1482\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1191\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1038\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_584\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1028\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_974\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1697\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1222_2\ : std_logic ;
  signal N_32777 : std_logic ;
  signal N_32980_1 : std_logic ;
  signal N_33734_1 : std_logic ;
  signal N_32904_2 : std_logic ;
  signal N_33140_1 : std_logic ;
  signal N_32844_2 : std_logic ;
  signal N_33219 : std_logic ;
  signal N_33253 : std_logic ;
  signal N_28652_1 : std_logic ;
  signal N_33427 : std_logic ;
  signal N_33368_1 : std_logic ;
  signal N_32727_1 : std_logic ;
  signal N_33431 : std_logic ;
  signal N_33504 : std_logic ;
  signal N_33510 : std_logic ;
  signal N_32908_1 : std_logic ;
  signal N_28211_1 : std_logic ;
  signal N_33507_1 : std_logic ;
  signal N_33647 : std_logic ;
  signal N_33733 : std_logic ;
  signal N_33833 : std_logic ;
  signal N_33899_1 : std_logic ;
  signal N_33902 : std_logic ;
  signal N_32738_1 : std_logic ;
  signal N_33968 : std_logic ;
  signal N_33074_1 : std_logic ;
  signal N_34263_2 : std_logic ;
  signal N_34040_1 : std_logic ;
  signal N_34043_2 : std_logic ;
  signal N_34257 : std_logic ;
  signal N_34325_1 : std_logic ;
  signal N_32861_1 : std_logic ;
  signal N_28251_1 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_531\ : std_logic ;
  signal N_34326_2 : std_logic ;
  signal N_33721_1 : std_logic ;
  signal N_28658_1 : std_logic ;
  signal N_34330 : std_logic ;
  signal N_34343_1 : std_logic ;
  signal N_34340_2 : std_logic ;
  signal N_34339_3 : std_logic ;
  signal N_34337 : std_logic ;
  signal N_34335_2 : std_logic ;
  signal N_28921_1 : std_logic ;
  signal N_34333 : std_logic ;
  signal N_32731_1 : std_logic ;
  signal N_32786_1 : std_logic ;
  signal N_34329 : std_logic ;
  signal N_34329_1 : std_logic ;
  signal N_34327 : std_logic ;
  signal N_34311_I : std_logic ;
  signal N_34279 : std_logic ;
  signal N_34272_1 : std_logic ;
  signal N_34271 : std_logic ;
  signal N_33070_1 : std_logic ;
  signal N_33718_1 : std_logic ;
  signal N_34268 : std_logic ;
  signal N_34262 : std_logic ;
  signal N_34260 : std_logic ;
  signal N_34259 : std_logic ;
  signal N_34239_I : std_logic ;
  signal N_34256_1 : std_logic ;
  signal N_34254 : std_logic ;
  signal N_34254_1 : std_logic ;
  signal N_34195 : std_logic ;
  signal N_34195_1 : std_logic ;
  signal N_34194 : std_logic ;
  signal N_34191 : std_logic ;
  signal N_33340_I : std_logic ;
  signal N_34190 : std_logic ;
  signal N_34187 : std_logic ;
  signal N_34184 : std_logic ;
  signal N_34183 : std_logic ;
  signal N_34182 : std_logic ;
  signal N_34181 : std_logic ;
  signal N_34180 : std_logic ;
  signal N_34133_2 : std_logic ;
  signal N_34132_1 : std_logic ;
  signal N_32791_1 : std_logic ;
  signal N_28250_2 : std_logic ;
  signal N_33447_1 : std_logic ;
  signal N_34029 : std_logic ;
  signal N_34127 : std_logic ;
  signal N_33735_1 : std_logic ;
  signal N_34123 : std_logic ;
  signal N_34121 : std_logic ;
  signal N_34120 : std_logic ;
  signal N_34119 : std_logic ;
  signal N_34118 : std_logic ;
  signal N_34117 : std_logic ;
  signal N_34114 : std_logic ;
  signal N_34113 : std_logic ;
  signal N_34111 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_719\ : std_logic ;
  signal N_34107 : std_logic ;
  signal N_34059 : std_logic ;
  signal N_34059_1 : std_logic ;
  signal N_34047_2 : std_logic ;
  signal N_34047 : std_logic ;
  signal N_34024 : std_logic ;
  signal N_34042 : std_logic ;
  signal N_34041 : std_logic ;
  signal N_34039 : std_logic ;
  signal N_33988_4 : std_logic ;
  signal N_28227_1 : std_logic ;
  signal N_33987 : std_logic ;
  signal N_33985_2 : std_logic ;
  signal N_33982 : std_logic ;
  signal N_34007 : std_logic ;
  signal N_33976 : std_logic ;
  signal N_33975 : std_logic ;
  signal N_33974 : std_logic ;
  signal N_32959_I : std_logic ;
  signal N_33973 : std_logic ;
  signal N_33972 : std_logic ;
  signal N_33971 : std_logic ;
  signal N_33970 : std_logic ;
  signal N_33967 : std_logic ;
  signal N_33966 : std_logic ;
  signal N_33914 : std_logic ;
  signal N_33913 : std_logic ;
  signal N_33668_1 : std_logic ;
  signal N_33912 : std_logic ;
  signal N_33911 : std_logic ;
  signal N_33870 : std_logic ;
  signal N_33908 : std_logic ;
  signal N_33905 : std_logic ;
  signal N_33900 : std_logic ;
  signal N_33897 : std_logic ;
  signal N_33896 : std_logic ;
  signal N_33503_1 : std_logic ;
  signal N_33895 : std_logic ;
  signal N_33847 : std_logic ;
  signal N_33845 : std_logic ;
  signal N_33844 : std_logic ;
  signal N_33842 : std_logic ;
  signal N_33841 : std_logic ;
  signal N_33839 : std_logic ;
  signal N_33838_2 : std_logic ;
  signal N_33834 : std_logic ;
  signal N_33832 : std_logic ;
  signal N_33830 : std_logic ;
  signal N_33813 : std_logic ;
  signal N_33828 : std_logic ;
  signal N_33827 : std_logic ;
  signal N_33777 : std_logic ;
  signal N_33795 : std_logic ;
  signal N_28681_I : std_logic ;
  signal N_32789_2 : std_logic ;
  signal N_33783 : std_logic ;
  signal N_33780 : std_logic ;
  signal N_33769 : std_logic ;
  signal N_33778 : std_logic ;
  signal N_33756 : std_logic ;
  signal N_33738_1 : std_logic ;
  signal N_33735_3 : std_logic ;
  signal N_33729 : std_logic ;
  signal N_33727_2 : std_logic ;
  signal N_33721 : std_logic ;
  signal N_33710 : std_logic ;
  signal N_33715 : std_logic ;
  signal N_33683 : std_logic ;
  signal N_33666 : std_logic ;
  signal N_33661 : std_logic ;
  signal N_33144_1 : std_logic ;
  signal N_33658 : std_logic ;
  signal N_33655 : std_logic ;
  signal N_33654 : std_logic ;
  signal N_33653 : std_logic ;
  signal N_33652 : std_logic ;
  signal N_33650 : std_logic ;
  signal N_33648 : std_logic ;
  signal N_33646 : std_logic ;
  signal N_33644 : std_logic ;
  signal N_33643 : std_logic ;
  signal N_28892_I : std_logic ;
  signal N_33590 : std_logic ;
  signal N_33589 : std_logic ;
  signal N_33588 : std_logic ;
  signal N_33584 : std_logic ;
  signal N_33547_I : std_logic ;
  signal N_33581 : std_logic ;
  signal N_33578 : std_logic ;
  signal N_33576 : std_logic ;
  signal N_33574 : std_logic ;
  signal N_33572 : std_logic ;
  signal N_33565 : std_logic ;
  signal N_33518 : std_logic ;
  signal N_33501_2 : std_logic ;
  signal N_33514 : std_logic ;
  signal N_33513 : std_logic ;
  signal N_33506 : std_logic ;
  signal N_33505 : std_logic ;
  signal N_33503 : std_logic ;
  signal N_33501 : std_logic ;
  signal N_33500 : std_logic ;
  signal N_33498 : std_logic ;
  signal N_33498_1 : std_logic ;
  signal N_33447 : std_logic ;
  signal N_33444 : std_logic ;
  signal N_28730_1 : std_logic ;
  signal N_33440 : std_logic ;
  signal N_33437 : std_logic ;
  signal N_33436 : std_logic ;
  signal N_33435 : std_logic ;
  signal N_33434 : std_logic ;
  signal N_33433 : std_logic ;
  signal N_33432 : std_logic ;
  signal N_33429 : std_logic ;
  signal N_33428 : std_logic ;
  signal N_33426 : std_logic ;
  signal N_33425 : std_logic ;
  signal N_33373 : std_logic ;
  signal N_33373_2 : std_logic ;
  signal N_33055 : std_logic ;
  signal N_33371 : std_logic ;
  signal N_33369 : std_logic ;
  signal N_33369_1 : std_logic ;
  signal N_33365 : std_logic ;
  signal N_33363 : std_logic ;
  signal N_33362 : std_logic ;
  signal N_33360 : std_logic ;
  signal N_33360_1 : std_logic ;
  signal N_33359 : std_logic ;
  signal N_33358 : std_logic ;
  signal N_33357 : std_logic ;
  signal N_33353 : std_logic ;
  signal N_33351 : std_logic ;
  signal N_33263_I : std_logic ;
  signal N_33297 : std_logic ;
  signal N_33293_2 : std_logic ;
  signal N_33291 : std_logic ;
  signal N_33289 : std_logic ;
  signal N_33288 : std_logic ;
  signal N_33286 : std_logic ;
  signal N_33277 : std_logic ;
  signal N_33283 : std_logic ;
  signal N_33278 : std_logic ;
  signal N_33229 : std_logic ;
  signal N_33225 : std_logic ;
  signal N_33224 : std_logic ;
  signal N_33220 : std_logic ;
  signal N_33217 : std_logic ;
  signal N_33215 : std_logic ;
  signal N_33210 : std_logic ;
  signal N_33209 : std_logic ;
  signal N_33208 : std_logic ;
  signal N_33149 : std_logic ;
  signal N_33148 : std_logic ;
  signal N_33125 : std_logic ;
  signal N_33123_1 : std_logic ;
  signal N_33081 : std_logic ;
  signal N_33079 : std_logic ;
  signal N_33076 : std_logic ;
  signal N_33073 : std_logic ;
  signal N_33071 : std_logic ;
  signal N_33070 : std_logic ;
  signal N_33069 : std_logic ;
  signal N_33068 : std_logic ;
  signal N_33061 : std_logic ;
  signal N_33022 : std_logic ;
  signal N_33032 : std_logic ;
  signal N_33031 : std_logic ;
  signal N_33028 : std_logic ;
  signal N_33027 : std_logic ;
  signal N_33026 : std_logic ;
  signal N_33024 : std_logic ;
  signal N_33021 : std_logic ;
  signal N_32982 : std_logic ;
  signal N_32981 : std_logic ;
  signal N_32981_1 : std_logic ;
  signal N_32976 : std_logic ;
  signal N_32956_I : std_logic ;
  signal N_32974 : std_logic ;
  signal N_32974_2 : std_logic ;
  signal N_32973 : std_logic ;
  signal N_32972 : std_logic ;
  signal N_32970 : std_logic ;
  signal N_32921 : std_logic ;
  signal N_32917 : std_logic ;
  signal N_32916 : std_logic ;
  signal N_32915 : std_logic ;
  signal N_32914 : std_logic ;
  signal N_32912 : std_logic ;
  signal N_32909 : std_logic ;
  signal N_32908 : std_logic ;
  signal N_32907 : std_logic ;
  signal N_32906 : std_logic ;
  signal N_32946 : std_logic ;
  signal N_32903 : std_logic ;
  signal N_32902 : std_logic ;
  signal N_32847 : std_logic ;
  signal N_32844 : std_logic ;
  signal N_32843 : std_logic ;
  signal N_32842 : std_logic ;
  signal N_32840_2 : std_logic ;
  signal N_32798 : std_logic ;
  signal N_32797 : std_logic ;
  signal N_32796_3 : std_logic ;
  signal N_32794 : std_logic ;
  signal N_32792 : std_logic ;
  signal N_32788 : std_logic ;
  signal N_32787 : std_logic ;
  signal N_32785 : std_logic ;
  signal N_32783 : std_logic ;
  signal N_32762_I : std_logic ;
  signal N_32780 : std_logic ;
  signal N_32735 : std_logic ;
  signal N_32732 : std_logic ;
  signal N_32732_2 : std_logic ;
  signal N_32731 : std_logic ;
  signal N_32729 : std_logic ;
  signal N_32727 : std_logic ;
  signal N_28207 : std_logic ;
  signal N_28206 : std_logic ;
  signal N_28212 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_571\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1048\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1714\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1049\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_467\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9375\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1592\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1082\ : std_logic ;
  signal N_28312_1 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1133\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1672\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1200\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1212\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1214\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1233\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1388\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1749\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1744\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_693\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1031\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1278\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1134\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9479\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1201\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_756\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1030\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1027\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8714\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1194\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_758\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8573\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_759\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1302\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1303\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1301\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1832\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1389\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8631\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9349\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9517\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1685\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_907\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1718\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9371\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11810_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9327\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8556\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9607\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9645\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9608\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9665\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8666\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9062\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9373\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8834\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8941\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9166\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9198\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9201\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8537\ : std_logic ;
  signal N_28212_1_0 : std_logic ;
  signal N_28242 : std_logic ;
  signal N_28251 : std_logic ;
  signal N_28252 : std_logic ;
  signal N_28253 : std_logic ;
  signal N_28254 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9368\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1682\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1595\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1568\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9511\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1800\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1206\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9547\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1135\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1054\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9099\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1234\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1236\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1235\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1036\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9397\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1079\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_948\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1053\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1044\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9157\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8619\ : std_logic ;
  signal N_33560 : std_logic ;
  signal N_28390_2 : std_logic ;
  signal N_28267 : std_logic ;
  signal N_28263 : std_logic ;
  signal N_28227 : std_logic ;
  signal N_28226 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_811\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_661\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1647\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1648\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1374\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1588\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_493\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1713\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1768\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9095_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1734\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9522\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9570\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9523\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7777\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7778\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7786\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10931\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_446\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_492\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10870\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10936\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TEMP\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.REEXCOVUV.UN25_LOCOV_0\ : std_logic ;
  signal \GRLFPC2_0.N_1391\ : std_logic ;
  signal \GRLFPC2_0.WREN2_2_SQMUXA\ : std_logic ;
  signal \GRLFPC2_0.N_1105\ : std_logic ;
  signal \GRLFPC2_0.N_71\ : std_logic ;
  signal \GRLFPC2_0.N_3091\ : std_logic ;
  signal \GRLFPC2_0.N_3423\ : std_logic ;
  signal \GRLFPC2_0.N_3097\ : std_logic ;
  signal \GRLFPC2_0.N_3099\ : std_logic ;
  signal \GRLFPC2_0.V.STATE_1_SQMUXA_3\ : std_logic ;
  signal \GRLFPC2_0.N_1667\ : std_logic ;
  signal \GRLFPC2_0.N_67\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9817\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9994\ : std_logic ;
  signal \GRLFPC2_0.N_82\ : std_logic ;
  signal N_37318_1 : std_logic ;
  signal \GRLFPC2_0.COMB.ISFPOP2_1\ : std_logic ;
  signal \GRLFPC2_0.N_1439\ : std_logic ;
  signal \GRLFPC2_0.N_1133\ : std_logic ;
  signal \GRLFPC2_0.N_58\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10503\ : std_logic ;
  signal \GRLFPC2_0.N_3077\ : std_logic ;
  signal \GRLFPC2_0.N_3106\ : std_logic ;
  signal \GRLFPC2_0.N_3093\ : std_logic ;
  signal \GRLFPC2_0.N_3429\ : std_logic ;
  signal \GRLFPC2_0.N_1495\ : std_logic ;
  signal N_37317 : std_logic ;
  signal \GRLFPC2_0.N_1438_15\ : std_logic ;
  signal \GRLFPC2_0.COMB.ANNULRES_1\ : std_logic ;
  signal \GRLFPC2_0.N_2888\ : std_logic ;
  signal \GRLFPC2_0.N_925\ : std_logic ;
  signal \GRLFPC2_0.N_43\ : std_logic ;
  signal \GRLFPC2_0.N_3466\ : std_logic ;
  signal \GRLFPC2_0.N_3468\ : std_logic ;
  signal \GRLFPC2_0.N_40\ : std_logic ;
  signal \GRLFPC2_0.N_44\ : std_logic ;
  signal \GRLFPC2_0.N_45\ : std_logic ;
  signal \GRLFPC2_0.COMB.RDD_1.N_27\ : std_logic ;
  signal \GRLFPC2_0.N_624_3\ : std_logic ;
  signal \GRLFPC2_0.RS1D_CNST\ : std_logic ;
  signal \GRLFPC2_0.COMB.RDD_1.N_12\ : std_logic ;
  signal \GRLFPC2_0.COMB.FPDECODE.RS1D5_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3924\ : std_logic ;
  signal N_37362 : std_logic ;
  signal \GRLFPC2_0.N_2975\ : std_logic ;
  signal N_37405 : std_logic ;
  signal N_37365_1 : std_logic ;
  signal \GRLFPC2_0.N_3462\ : std_logic ;
  signal \GRLFPC2_0.RS1V_0_SQMUXA\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_959_I\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN26_GEN\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5452\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5458\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5771\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6583\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP_1_1_CO1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5446\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1618\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10902\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10909\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_663\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10881\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1493\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_429\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1495\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1497\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1637\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1509\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1636\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1844\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1633\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_504\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1677\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1770\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1771\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1836\ : std_logic ;
  signal N_35132 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_547\ : std_logic ;
  signal N_28511 : std_logic ;
  signal N_28510 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1505\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_451\ : std_logic ;
  signal N_35133 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1496\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1492\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1515\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1516\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1518\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1519\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1520\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1503\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1839\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1852\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1544\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1846\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_743\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_386\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_389\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_893\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10879\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10864\ : std_logic ;
  signal \GRLFPC2_0.N_1714_I\ : std_logic ;
  signal \GRLFPC2_0.N_1093\ : std_logic ;
  signal \GRLFPC2_0.N_1072\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1855\ : std_logic ;
  signal \GRLFPC2_0.N_3475\ : std_logic ;
  signal \GRLFPC2_0.N_3027\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_1\ : std_logic ;
  signal \GRLFPC2_0.FPI.RST_1\ : std_logic ;
  signal \GRLFPC2_0.R.MK.RST_4\ : std_logic ;
  signal \GRLFPC2_0.N_3545\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5335\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10882\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3639\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10525\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10527\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6961\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10626\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN11_WQSTSETS\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4534\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_1_CO0\ : std_logic ;
  signal \GRLFPC2_0.N_77_1\ : std_logic ;
  signal N_37387 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4662\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5343\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5339\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5301\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC\ : std_logic ;
  signal \GRLFPC2_0.V.FSR.CEXC_2_SQMUXA\ : std_logic ;
  signal N_37320 : std_logic ;
  signal \GRLFPC2_0.R.I.V_1_0_G2\ : std_logic ;
  signal \GRLFPC2_0.V.FSR.CEXC_3_SQMUXA\ : std_logic ;
  signal \GRLFPC2_0.N_3114\ : std_logic ;
  signal \GRLFPC2_0.N_3432\ : std_logic ;
  signal \GRLFPC2_0.N_3052\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10523\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10522\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10524\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10521\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10520\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10519\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10518\ : std_logic ;
  signal \GRLFPC2_0.N_3086\ : std_logic ;
  signal \GRLFPC2_0.N_3054\ : std_logic ;
  signal \GRLFPC2_0.N_3433\ : std_logic ;
  signal \GRLFPC2_0.N_3056\ : std_logic ;
  signal \GRLFPC2_0.N_3090\ : std_logic ;
  signal \GRLFPC2_0.N_3059\ : std_logic ;
  signal \GRLFPC2_0.N_3434\ : std_logic ;
  signal \GRLFPC2_0.N_3435\ : std_logic ;
  signal \GRLFPC2_0.N_3436\ : std_logic ;
  signal \GRLFPC2_0.N_3437\ : std_logic ;
  signal \GRLFPC2_0.N_3439\ : std_logic ;
  signal \GRLFPC2_0.N_3101\ : std_logic ;
  signal \GRLFPC2_0.N_3069\ : std_logic ;
  signal \GRLFPC2_0.N_3103\ : std_logic ;
  signal \GRLFPC2_0.N_3442\ : std_logic ;
  signal \GRLFPC2_0.N_3443\ : std_logic ;
  signal \GRLFPC2_0.N_3445\ : std_logic ;
  signal \GRLFPC2_0.N_3108\ : std_logic ;
  signal \GRLFPC2_0.N_3109\ : std_logic ;
  signal \GRLFPC2_0.N_3078\ : std_logic ;
  signal \GRLFPC2_0.N_3079\ : std_logic ;
  signal \GRLFPC2_0.N_3446\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897\ : std_logic ;
  signal \GRLFPC2_0.N_3227\ : std_logic ;
  signal \GRLFPC2_0.N_3426\ : std_logic ;
  signal \GRLFPC2_0.N_3425\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN31_DEBUG_UNIT\ : std_logic ;
  signal \GRLFPC2_0.N_3226\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10006\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9991\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9820\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9997\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9963\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9822\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10206\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9968\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9962\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9961\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9979\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9973\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9972\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9984\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9982\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9990\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10005\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10002\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9999\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9995\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9992\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9977\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10001\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10008\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9975\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9978\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10204\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10203\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9966\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9960\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9971\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9974\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9985\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10010\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10195\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9782\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9781\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10207\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9789\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9980\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9805\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10009\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10878\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10877\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10880\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10514\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10512\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10197\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9783\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10004\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9967\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10003\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9986\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9970\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9987\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10000\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9976\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9964\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9988\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10007\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10934\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10862\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10876\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10875\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10861\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10874\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10860\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10873\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10857\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10011\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9989\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9983\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10859\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10872\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10858\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10871\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9969\ : std_logic ;
  signal \GRLFPC2_0.FPO.SIGN\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_60.Z_1_CO1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1281_I\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7035\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_402\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1539\ : std_logic ;
  signal \GRLFPC2_0.N_74\ : std_logic ;
  signal \GRLFPC2_0.N_94\ : std_logic ;
  signal \GRLFPC2_0.N_3458\ : std_logic ;
  signal \GRLFPC2_0.N_3491\ : std_logic ;
  signal \GRLFPC2_0.N_552_1_0\ : std_logic ;
  signal \GRLFPC2_0.N_1841\ : std_logic ;
  signal \GRLFPC2_0.N_90\ : std_logic ;
  signal \GRLFPC2_0.N_138\ : std_logic ;
  signal \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1540\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_875\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_403\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4664\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5416\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN40_SHDVAR\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN20_SHDVAR\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal N_30731 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1274_I\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4238\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN5_SHDVAR\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7051\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7034\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_12231\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN13_RESVEC\ : std_logic ;
  signal N_42365 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_TZ\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_4_TZ\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_1\ : std_logic ;
  signal N_44753 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S\ : std_logic ;
  signal N_44786 : std_logic ;
  signal N_44787 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3\ : std_logic ;
  signal D_N_7 : std_logic ;
  signal \GRLFPC2_0.RS1V12_TZ\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_5_TZ\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_6_TZ\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_8_TZ\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_4_TZ\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_11_TZ\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_18_TZ\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0_N_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_13_TZ\ : std_logic ;
  signal \GRLFPC2_0.WREN2_1_SQMUXA_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.A.RF2REN_1_8055_I_A5_0_0\ : std_logic ;
  signal N_33725_1 : std_logic ;
  signal N_33652_1 : std_logic ;
  signal N_33222_2 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9490\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9492\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.STATE12_0\ : std_logic ;
  signal N_37019_2 : std_logic ;
  signal N_52053 : std_logic ;
  signal N_52054 : std_logic ;
  signal N_52055 : std_logic ;
  signal N_52056 : std_logic ;
  signal N_52057 : std_logic ;
  signal N_52058 : std_logic ;
  signal N_52059 : std_logic ;
  signal N_52060 : std_logic ;
  signal N_52061 : std_logic ;
  signal N_52062 : std_logic ;
  signal N_52063 : std_logic ;
  signal N_52064 : std_logic ;
  signal N_52065 : std_logic ;
  signal N_52066 : std_logic ;
  signal N_52067 : std_logic ;
  signal N_52068 : std_logic ;
  signal N_52069 : std_logic ;
  signal N_52070 : std_logic ;
  signal N_52071 : std_logic ;
  signal N_52072 : std_logic ;
  signal N_52073 : std_logic ;
  signal N_52074 : std_logic ;
  signal N_52075 : std_logic ;
  signal N_52076 : std_logic ;
  signal N_52079 : std_logic ;
  signal N_52080 : std_logic ;
  signal N_52081 : std_logic ;
  signal N_52082 : std_logic ;
  signal N_52083 : std_logic ;
  signal N_52084 : std_logic ;
  signal N_52085 : std_logic ;
  signal N_52086 : std_logic ;
  signal N_52087 : std_logic ;
  signal N_52088 : std_logic ;
  signal N_52089 : std_logic ;
  signal N_52090 : std_logic ;
  signal N_52091 : std_logic ;
  signal N_52092 : std_logic ;
  signal N_52093 : std_logic ;
  signal N_52094 : std_logic ;
  signal N_52095 : std_logic ;
  signal N_52096 : std_logic ;
  signal N_52097 : std_logic ;
  signal N_52098 : std_logic ;
  signal N_52099 : std_logic ;
  signal N_52100 : std_logic ;
  signal N_52101 : std_logic ;
  signal N_52102 : std_logic ;
  signal N_52103 : std_logic ;
  signal N_52104 : std_logic ;
  signal N_52105 : std_logic ;
  signal N_52106 : std_logic ;
  signal N_52107 : std_logic ;
  signal N_52108 : std_logic ;
  signal N_52109 : std_logic ;
  signal N_52110 : std_logic ;
  signal N_52111 : std_logic ;
  signal N_52112 : std_logic ;
  signal N_52113 : std_logic ;
  signal N_52114 : std_logic ;
  signal N_52115 : std_logic ;
  signal N_52116 : std_logic ;
  signal N_52117 : std_logic ;
  signal N_52118 : std_logic ;
  signal N_52119 : std_logic ;
  signal N_52120 : std_logic ;
  signal N_52121 : std_logic ;
  signal N_52122 : std_logic ;
  signal N_52123 : std_logic ;
  signal N_52124 : std_logic ;
  signal N_52125 : std_logic ;
  signal N_52126 : std_logic ;
  signal N_52127 : std_logic ;
  signal N_52128 : std_logic ;
  signal N_52129 : std_logic ;
  signal N_52130 : std_logic ;
  signal N_52131 : std_logic ;
  signal N_52132 : std_logic ;
  signal N_52133 : std_logic ;
  signal N_52134 : std_logic ;
  signal N_52135 : std_logic ;
  signal N_52136 : std_logic ;
  signal N_52137 : std_logic ;
  signal N_52138 : std_logic ;
  signal N_52139 : std_logic ;
  signal N_52140 : std_logic ;
  signal N_52141 : std_logic ;
  signal N_52142 : std_logic ;
  signal N_52143 : std_logic ;
  signal N_52144 : std_logic ;
  signal N_52145 : std_logic ;
  signal N_52146 : std_logic ;
  signal N_52147 : std_logic ;
  signal N_52148 : std_logic ;
  signal N_52149 : std_logic ;
  signal N_52150 : std_logic ;
  signal N_52151 : std_logic ;
  signal N_52152 : std_logic ;
  signal N_52153 : std_logic ;
  signal N_52154 : std_logic ;
  signal N_52155 : std_logic ;
  signal N_52156 : std_logic ;
  signal N_52157 : std_logic ;
  signal N_52158 : std_logic ;
  signal N_52159 : std_logic ;
  signal N_52160 : std_logic ;
  signal N_52161 : std_logic ;
  signal N_52162 : std_logic ;
  signal N_52163 : std_logic ;
  signal N_52164 : std_logic ;
  signal N_52165 : std_logic ;
  signal N_52166 : std_logic ;
  signal N_52167 : std_logic ;
  signal N_52168 : std_logic ;
  signal N_52169 : std_logic ;
  signal N_52170 : std_logic ;
  signal N_52171 : std_logic ;
  signal N_52172 : std_logic ;
  signal N_52173 : std_logic ;
  signal N_52174 : std_logic ;
  signal N_52175 : std_logic ;
  signal N_52176 : std_logic ;
  signal N_52177 : std_logic ;
  signal N_52178 : std_logic ;
  signal N_52179 : std_logic ;
  signal N_52180 : std_logic ;
  signal N_52181 : std_logic ;
  signal N_52182 : std_logic ;
  signal N_52183 : std_logic ;
  signal N_52184 : std_logic ;
  signal N_52185 : std_logic ;
  signal N_52186 : std_logic ;
  signal N_52187 : std_logic ;
  signal N_52188 : std_logic ;
  signal N_52189 : std_logic ;
  signal N_52190 : std_logic ;
  signal N_52191 : std_logic ;
  signal N_52192 : std_logic ;
  signal N_52193 : std_logic ;
  signal N_52194 : std_logic ;
  signal N_52195 : std_logic ;
  signal N_52196 : std_logic ;
  signal N_52197 : std_logic ;
  signal N_52198 : std_logic ;
  signal N_52199 : std_logic ;
  signal N_52200 : std_logic ;
  signal N_52201 : std_logic ;
  signal N_52202 : std_logic ;
  signal N_52203 : std_logic ;
  signal N_52204 : std_logic ;
  signal N_52205 : std_logic ;
  signal N_52206 : std_logic ;
  signal N_52207 : std_logic ;
  signal N_52208 : std_logic ;
  signal N_52209 : std_logic ;
  signal N_52210 : std_logic ;
  signal N_52211 : std_logic ;
  signal N_52212 : std_logic ;
  signal N_52213 : std_logic ;
  signal N_52214 : std_logic ;
  signal N_52215 : std_logic ;
  signal N_52216 : std_logic ;
  signal N_52217 : std_logic ;
  signal N_52218 : std_logic ;
  signal N_52219 : std_logic ;
  signal N_52220 : std_logic ;
  signal N_52221 : std_logic ;
  signal N_52222 : std_logic ;
  signal N_52223 : std_logic ;
  signal N_52224 : std_logic ;
  signal N_52225 : std_logic ;
  signal N_52226 : std_logic ;
  signal N_52227 : std_logic ;
  signal N_52228 : std_logic ;
  signal N_52229 : std_logic ;
  signal N_52230 : std_logic ;
  signal N_52231 : std_logic ;
  signal N_52232 : std_logic ;
  signal N_52233 : std_logic ;
  signal N_52234 : std_logic ;
  signal N_52235 : std_logic ;
  signal N_52236 : std_logic ;
  signal N_52237 : std_logic ;
  signal N_52238 : std_logic ;
  signal N_52239 : std_logic ;
  signal N_52240 : std_logic ;
  signal N_52241 : std_logic ;
  signal N_52242 : std_logic ;
  signal N_52243 : std_logic ;
  signal N_52244 : std_logic ;
  signal N_52245 : std_logic ;
  signal N_52246 : std_logic ;
  signal N_52247 : std_logic ;
  signal N_52248 : std_logic ;
  signal N_52249 : std_logic ;
  signal N_52250 : std_logic ;
  signal N_52251 : std_logic ;
  signal N_52252 : std_logic ;
  signal N_52253 : std_logic ;
  signal N_52254 : std_logic ;
  signal N_52255 : std_logic ;
  signal N_52256 : std_logic ;
  signal N_52257 : std_logic ;
  signal N_52258 : std_logic ;
  signal N_52259 : std_logic ;
  signal N_52260 : std_logic ;
  signal N_52261 : std_logic ;
  signal N_52262 : std_logic ;
  signal N_52263 : std_logic ;
  signal N_52264 : std_logic ;
  signal N_52265 : std_logic ;
  signal N_52266 : std_logic ;
  signal N_52267 : std_logic ;
  signal N_52268 : std_logic ;
  signal N_52272 : std_logic ;
  signal N_52273 : std_logic ;
  signal N_52279 : std_logic ;
  signal N_52280 : std_logic ;
  signal N_52288 : std_logic ;
  signal N_52295 : std_logic ;
  signal N_52296 : std_logic ;
  signal N_52302 : std_logic ;
  signal N_52303 : std_logic ;
  signal N_52311 : std_logic ;
  signal N_52318 : std_logic ;
  signal N_52319 : std_logic ;
  signal N_52325 : std_logic ;
  signal N_52326 : std_logic ;
  signal N_52334 : std_logic ;
  signal N_52341 : std_logic ;
  signal N_52342 : std_logic ;
  signal N_52348 : std_logic ;
  signal N_52349 : std_logic ;
  signal N_52357 : std_logic ;
  signal N_52364 : std_logic ;
  signal N_52365 : std_logic ;
  signal N_52371 : std_logic ;
  signal N_52372 : std_logic ;
  signal N_52380 : std_logic ;
  signal N_52387 : std_logic ;
  signal N_52388 : std_logic ;
  signal N_52394 : std_logic ;
  signal N_52395 : std_logic ;
  signal N_52403 : std_logic ;
  signal N_52410 : std_logic ;
  signal N_52411 : std_logic ;
  signal N_52417 : std_logic ;
  signal N_52418 : std_logic ;
  signal N_52426 : std_logic ;
  signal N_52433 : std_logic ;
  signal N_52434 : std_logic ;
  signal N_52440 : std_logic ;
  signal N_52441 : std_logic ;
  signal N_52449 : std_logic ;
  signal N_52456 : std_logic ;
  signal N_52457 : std_logic ;
  signal N_52463 : std_logic ;
  signal N_52464 : std_logic ;
  signal N_52472 : std_logic ;
  signal N_52479 : std_logic ;
  signal N_52480 : std_logic ;
  signal N_52486 : std_logic ;
  signal N_52487 : std_logic ;
  signal N_52495 : std_logic ;
  signal N_52502 : std_logic ;
  signal N_52503 : std_logic ;
  signal N_52509 : std_logic ;
  signal N_52510 : std_logic ;
  signal N_52518 : std_logic ;
  signal N_52525 : std_logic ;
  signal N_52526 : std_logic ;
  signal N_52532 : std_logic ;
  signal N_52533 : std_logic ;
  signal N_52541 : std_logic ;
  signal N_52548 : std_logic ;
  signal N_52549 : std_logic ;
  signal N_52555 : std_logic ;
  signal N_52556 : std_logic ;
  signal N_52564 : std_logic ;
  signal N_52571 : std_logic ;
  signal N_52572 : std_logic ;
  signal N_52578 : std_logic ;
  signal N_52579 : std_logic ;
  signal N_52587 : std_logic ;
  signal N_52594 : std_logic ;
  signal N_52595 : std_logic ;
  signal N_52601 : std_logic ;
  signal N_52602 : std_logic ;
  signal N_52610 : std_logic ;
  signal N_52617 : std_logic ;
  signal N_52618 : std_logic ;
  signal N_52624 : std_logic ;
  signal N_52625 : std_logic ;
  signal N_52633 : std_logic ;
  signal N_52640 : std_logic ;
  signal N_52641 : std_logic ;
  signal N_52647 : std_logic ;
  signal N_52648 : std_logic ;
  signal N_52656 : std_logic ;
  signal N_52663 : std_logic ;
  signal N_52664 : std_logic ;
  signal N_52670 : std_logic ;
  signal N_52671 : std_logic ;
  signal N_52679 : std_logic ;
  signal N_52686 : std_logic ;
  signal N_52687 : std_logic ;
  signal N_52693 : std_logic ;
  signal N_52694 : std_logic ;
  signal N_52702 : std_logic ;
  signal N_52709 : std_logic ;
  signal N_52710 : std_logic ;
  signal N_52716 : std_logic ;
  signal N_52717 : std_logic ;
  signal N_52725 : std_logic ;
  signal N_52732 : std_logic ;
  signal N_52733 : std_logic ;
  signal N_52739 : std_logic ;
  signal N_52740 : std_logic ;
  signal N_52748 : std_logic ;
  signal N_52755 : std_logic ;
  signal N_52756 : std_logic ;
  signal N_52762 : std_logic ;
  signal N_52763 : std_logic ;
  signal N_52771 : std_logic ;
  signal N_52778 : std_logic ;
  signal N_52779 : std_logic ;
  signal N_52785 : std_logic ;
  signal N_52786 : std_logic ;
  signal N_52794 : std_logic ;
  signal N_52801 : std_logic ;
  signal N_52802 : std_logic ;
  signal N_52808 : std_logic ;
  signal N_52809 : std_logic ;
  signal N_52817 : std_logic ;
  signal N_52824 : std_logic ;
  signal N_52825 : std_logic ;
  signal N_52831 : std_logic ;
  signal N_52832 : std_logic ;
  signal N_52840 : std_logic ;
  signal N_52847 : std_logic ;
  signal N_52848 : std_logic ;
  signal N_52854 : std_logic ;
  signal N_52855 : std_logic ;
  signal N_52863 : std_logic ;
  signal N_52870 : std_logic ;
  signal N_52871 : std_logic ;
  signal N_52877 : std_logic ;
  signal N_52878 : std_logic ;
  signal N_52886 : std_logic ;
  signal N_52893 : std_logic ;
  signal N_52894 : std_logic ;
  signal N_52900 : std_logic ;
  signal N_52901 : std_logic ;
  signal N_52909 : std_logic ;
  signal N_52916 : std_logic ;
  signal N_52917 : std_logic ;
  signal N_52923 : std_logic ;
  signal N_52924 : std_logic ;
  signal N_52932 : std_logic ;
  signal N_52939 : std_logic ;
  signal N_52940 : std_logic ;
  signal N_52946 : std_logic ;
  signal N_52947 : std_logic ;
  signal N_52955 : std_logic ;
  signal N_52962 : std_logic ;
  signal N_52963 : std_logic ;
  signal N_52969 : std_logic ;
  signal N_52970 : std_logic ;
  signal N_52978 : std_logic ;
  signal N_52985 : std_logic ;
  signal N_52986 : std_logic ;
  signal N_52992 : std_logic ;
  signal N_52993 : std_logic ;
  signal N_53001 : std_logic ;
  signal N_53008 : std_logic ;
  signal N_53009 : std_logic ;
  signal N_53015 : std_logic ;
  signal N_53016 : std_logic ;
  signal N_53024 : std_logic ;
  signal N_53034 : std_logic ;
  signal N_53044 : std_logic ;
  signal N_53045 : std_logic ;
  signal N_53048 : std_logic ;
  signal N_53049 : std_logic ;
  signal N_53053 : std_logic ;
  signal N_53054 : std_logic ;
  signal N_53060 : std_logic ;
  signal N_53061 : std_logic ;
  signal N_53069 : std_logic ;
  signal N_53076 : std_logic ;
  signal N_53077 : std_logic ;
  signal N_53083 : std_logic ;
  signal N_53084 : std_logic ;
  signal N_53092 : std_logic ;
  signal N_53099 : std_logic ;
  signal N_53100 : std_logic ;
  signal N_53106 : std_logic ;
  signal N_53107 : std_logic ;
  signal N_53115 : std_logic ;
  signal N_53122 : std_logic ;
  signal N_53123 : std_logic ;
  signal N_53129 : std_logic ;
  signal N_53130 : std_logic ;
  signal N_53138 : std_logic ;
  signal N_53145 : std_logic ;
  signal N_53146 : std_logic ;
  signal N_53152 : std_logic ;
  signal N_53153 : std_logic ;
  signal N_53161 : std_logic ;
  signal N_53168 : std_logic ;
  signal N_53169 : std_logic ;
  signal N_53175 : std_logic ;
  signal N_53176 : std_logic ;
  signal N_53184 : std_logic ;
  signal N_53191 : std_logic ;
  signal N_53192 : std_logic ;
  signal N_53198 : std_logic ;
  signal N_53199 : std_logic ;
  signal N_53207 : std_logic ;
  signal N_53214 : std_logic ;
  signal N_53215 : std_logic ;
  signal N_53221 : std_logic ;
  signal N_53222 : std_logic ;
  signal N_53230 : std_logic ;
  signal N_53237 : std_logic ;
  signal N_53238 : std_logic ;
  signal N_53244 : std_logic ;
  signal N_53245 : std_logic ;
  signal N_53253 : std_logic ;
  signal N_53260 : std_logic ;
  signal N_53261 : std_logic ;
  signal N_53267 : std_logic ;
  signal N_53268 : std_logic ;
  signal N_53276 : std_logic ;
  signal N_53283 : std_logic ;
  signal N_53284 : std_logic ;
  signal N_53290 : std_logic ;
  signal N_53291 : std_logic ;
  signal N_53299 : std_logic ;
  signal N_53306 : std_logic ;
  signal N_53307 : std_logic ;
  signal N_53313 : std_logic ;
  signal N_53314 : std_logic ;
  signal N_53322 : std_logic ;
  signal N_53329 : std_logic ;
  signal N_53330 : std_logic ;
  signal N_53336 : std_logic ;
  signal N_53337 : std_logic ;
  signal N_53345 : std_logic ;
  signal N_53416 : std_logic ;
  signal N_53417 : std_logic ;
  signal N_53423 : std_logic ;
  signal N_53424 : std_logic ;
  signal N_53434 : std_logic ;
  signal N_53435 : std_logic ;
  signal N_53441 : std_logic ;
  signal N_53442 : std_logic ;
  signal N_53450 : std_logic ;
  signal N_53457 : std_logic ;
  signal N_53458 : std_logic ;
  signal N_53464 : std_logic ;
  signal N_53465 : std_logic ;
  signal N_53473 : std_logic ;
  signal N_53480 : std_logic ;
  signal N_53481 : std_logic ;
  signal N_53487 : std_logic ;
  signal N_53488 : std_logic ;
  signal N_53496 : std_logic ;
  signal N_53503 : std_logic ;
  signal N_53504 : std_logic ;
  signal N_53510 : std_logic ;
  signal N_53511 : std_logic ;
  signal N_53519 : std_logic ;
  signal N_53526 : std_logic ;
  signal N_53527 : std_logic ;
  signal N_53533 : std_logic ;
  signal N_53534 : std_logic ;
  signal N_53542 : std_logic ;
  signal N_37343_I_0 : std_logic ;
  signal \GRLFPC2_0.N_3477_1_I\ : std_logic ;
  signal CPI_D_INST_INTERNAL_6 : std_logic ;
  signal \GRLFPC2_0.N_1830_O\ : std_logic ;
  signal \GRLFPC2_0.N_1683\ : std_logic ;
  signal \GRLFPC2_0.N_1685\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7226\ : std_logic ;
  signal N_53873 : std_logic ;
  signal N_53874 : std_logic ;
  signal N_53875 : std_logic ;
  signal N_53877 : std_logic ;
  signal N_53878 : std_logic ;
  signal N_53879 : std_logic ;
  signal N_53880 : std_logic ;
  signal N_53882 : std_logic ;
  signal N_53883 : std_logic ;
  signal N_53884 : std_logic ;
  signal N_53885 : std_logic ;
  signal N_53886 : std_logic ;
  signal N_53887 : std_logic ;
  signal N_53888 : std_logic ;
  signal N_53889 : std_logic ;
  signal N_53890 : std_logic ;
  signal N_53891 : std_logic ;
  signal N_53892 : std_logic ;
  signal N_53895 : std_logic ;
  signal N_53896 : std_logic ;
  signal N_53898 : std_logic ;
  signal N_53901 : std_logic ;
  signal N_53903 : std_logic ;
  signal N_53904 : std_logic ;
  signal N_53905 : std_logic ;
  signal N_53907 : std_logic ;
  signal N_53908 : std_logic ;
  signal N_53909 : std_logic ;
  signal N_53911 : std_logic ;
  signal N_53912 : std_logic ;
  signal N_53913 : std_logic ;
  signal N_53914 : std_logic ;
  signal N_53915 : std_logic ;
  signal N_53916 : std_logic ;
  signal N_53917 : std_logic ;
  signal N_53919 : std_logic ;
  signal N_53922 : std_logic ;
  signal N_53923 : std_logic ;
  signal N_53924 : std_logic ;
  signal N_53925 : std_logic ;
  signal N_53926 : std_logic ;
  signal N_53927 : std_logic ;
  signal N_53929 : std_logic ;
  signal N_53930 : std_logic ;
  signal N_53931 : std_logic ;
  signal N_53932 : std_logic ;
  signal N_53933 : std_logic ;
  signal N_53935 : std_logic ;
  signal N_53938 : std_logic ;
  signal N_53942 : std_logic ;
  signal N_53945 : std_logic ;
  signal N_53946 : std_logic ;
  signal N_53947 : std_logic ;
  signal N_53948 : std_logic ;
  signal N_53952 : std_logic ;
  signal N_53953 : std_logic ;
  signal N_53955 : std_logic ;
  signal N_53956 : std_logic ;
  signal N_53957 : std_logic ;
  signal N_53958 : std_logic ;
  signal N_53959 : std_logic ;
  signal N_53961 : std_logic ;
  signal N_53962 : std_logic ;
  signal N_53963 : std_logic ;
  signal N_53964 : std_logic ;
  signal N_53966 : std_logic ;
  signal N_53969 : std_logic ;
  signal N_53970 : std_logic ;
  signal N_53971 : std_logic ;
  signal N_53972 : std_logic ;
  signal N_53973 : std_logic ;
  signal N_53974 : std_logic ;
  signal N_53976 : std_logic ;
  signal N_53977 : std_logic ;
  signal N_53978 : std_logic ;
  signal N_53979 : std_logic ;
  signal N_53980 : std_logic ;
  signal N_53981 : std_logic ;
  signal N_53982 : std_logic ;
  signal N_53984 : std_logic ;
  signal N_53985 : std_logic ;
  signal N_53986 : std_logic ;
  signal N_53988 : std_logic ;
  signal N_53989 : std_logic ;
  signal N_53994 : std_logic ;
  signal N_53995 : std_logic ;
  signal N_53996 : std_logic ;
  signal N_53997 : std_logic ;
  signal N_53998 : std_logic ;
  signal N_53999 : std_logic ;
  signal N_54000 : std_logic ;
  signal N_54001 : std_logic ;
  signal N_54002 : std_logic ;
  signal N_54005 : std_logic ;
  signal N_54012 : std_logic ;
  signal N_54013 : std_logic ;
  signal N_54015 : std_logic ;
  signal N_54017 : std_logic ;
  signal N_54021 : std_logic ;
  signal N_54022 : std_logic ;
  signal N_54028 : std_logic ;
  signal N_54031 : std_logic ;
  signal N_54033 : std_logic ;
  signal N_54039 : std_logic ;
  signal N_54041 : std_logic ;
  signal N_54042 : std_logic ;
  signal N_54046 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_16_TZ\ : std_logic ;
  signal N_58999 : std_logic ;
  signal N_59000 : std_logic ;
  signal N_59001 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_10_TZ\ : std_logic ;
  signal \GRLFPC2_0.COMB.WREN1_9_IV_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.WREN1_9_IV_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.RDD_1.M7_E_54_I_A2_0_3\ : std_logic ;
  signal \GRLFPC2_0.UN1_FPOP7_1_0_A2_0_2\ : std_logic ;
  signal \GRLFPC2_0.COMB.WREN2_9_IV_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.WREN2_9_IV_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.RDD_1.M7_E_54_I_A2_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.A.RF1REN_1_8000_I_A5_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.FPDECODE.RS1D5_0_A2_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.RDD_1.M7_E_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN1_MEXC_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN1_MEXC_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7920_I_A7_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7920_I_A7_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7920_I_A7_10\ : std_logic ;
  signal \GRLFPC2_0.COMB.ANNULFPU_1_U_0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.I.RDD_1_I_A3_15_5_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.I.RDD_1_I_A3_15_7\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.I.RDD_1_I_A3_15_8\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.I.RDD_1_I_A3_15_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_19\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_20\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_22\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_23\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_26\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_27\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_28\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7920_I_1_1\ : std_logic ;
  signal \GRLFPC2_0.N_202\ : std_logic ;
  signal \GRLFPC2_0.R.E.AFQ_RET_0_0_G1_3\ : std_logic ;
  signal \GRLFPC2_0.R.E.AFQ_RET_0_0_G1_5\ : std_logic ;
  signal \GRLFPC2_0.R.A.LD_0_0_G1_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3945_I_I_O2_3_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN12_SRTOSTICKY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_14__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_24__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_39__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_44__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_19\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_18\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_19\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_13_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_16\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_16_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_18\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_20\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_22\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_18\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_18\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_20\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_18\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_11_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_16\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_18\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_11_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_15__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_6_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_8_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_19\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_13_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_18_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_20\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_21\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_23\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_30__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_30__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_10_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_16__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_16\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_17\ : std_logic ;
  signal \GRLFPC2_0.R.I.EXEC_0_0_G1_0_7945_I_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_8_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_16\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_20\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_22\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1_0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_12\ : std_logic ;
  signal \GRLFPC2_0.R.I.V_1_0_G0_I_O4_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_A2_7_8923_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_16\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_20\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_24\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_28\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_33\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_40\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_42\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_44\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_46\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_47\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_48\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_50\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_51\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_53\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__G2_0_7550_I_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_243__G2_0_7581_I_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_242__G2_0_7612_I_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_241__G2_0_7643_I_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_240__G2_0_7674_I_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.MIFROMINST_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_239__G2_0_7705_I_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_238__G2_0_7736_I_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_237__G2_0_7767_I_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_TZ_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.REEXCOVUV.UN13_LOCOV_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.REEXCOVUV.UN13_LOCOV_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN36_STKGEN_0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0_M3_I_A3_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_0_0_13__G0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.BUSYMULXFF.UN2_TEMP_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP\ : std_logic ;
  signal \GRLFPC2_0.N_1438\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5346\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN1_FPCI_4\ : std_logic ;
  signal \GRLFPC2_0.V.FSR.CEXC_0_SQMUXA\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\ : std_logic ;
  signal \GRLFPC2_0.N_951\ : std_logic ;
  signal \GRLFPC2_0.N_1243\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10530\ : std_logic ;
  signal \GRLFPC2_0.N_1171\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\ : std_logic ;
  signal \GRLFPC2_0.N_1517\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN1_R.A.RS1_1\ : std_logic ;
  signal \GRLFPC2_0.WRADDR_1_SQMUXA\ : std_logic ;
  signal \GRLFPC2_0.WRADDR_0_SQMUXA_1\ : std_logic ;
  signal \GRLFPC2_0.N_91\ : std_logic ;
  signal \GRLFPC2_0.N_1015\ : std_logic ;
  signal \GRLFPC2_0.N_83\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7352\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7350\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1586\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9525\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9486\ : std_logic ;
  signal N_33794 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_525\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9600\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9498\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\ : std_logic ;
  signal \GRLFPC2_0.N_1876_2\ : std_logic ;
  signal N_61580 : std_logic ;
  signal \GRLFPC2_0.R.I.INST_1_0_9__G2\ : std_logic ;
  signal \GRLFPC2_0.R.A.AFQ\ : std_logic ;
  signal \GRLFPC2_0.R.A.AFSR\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_473\ : std_logic ;
  signal N_61587_I : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\ : std_logic ;
  signal \GRLFPC2_0.N_54\ : std_logic ;
  signal N_65488 : std_logic ;
  signal N_65496 : std_logic ;
  signal N_65516 : std_logic ;
  signal N_65522 : std_logic ;
  signal N_65526 : std_logic ;
  signal N_65528 : std_logic ;
  signal N_65541 : std_logic ;
  signal N_65549 : std_logic ;
  signal N_65570 : std_logic ;
  signal N_65572 : std_logic ;
  signal N_65578 : std_logic ;
  signal N_65584 : std_logic ;
  signal N_65588 : std_logic ;
  signal N_65602 : std_logic ;
  signal N_65607 : std_logic ;
  signal N_65608 : std_logic ;
  signal N_65610 : std_logic ;
  signal N_65611 : std_logic ;
  signal N_65612 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6\ : std_logic ;
  signal N_65677 : std_logic ;
  signal N_65701 : std_logic ;
  signal N_65705 : std_logic ;
  signal N_65707 : std_logic ;
  signal N_65709 : std_logic ;
  signal N_65719 : std_logic ;
  signal N_65775 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_N_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_N_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10744\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10746\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10546\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10545\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7352_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO\ : std_logic ;
  signal N_1_0 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO\ : std_logic ;
  signal N_1_1 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO\ : std_logic ;
  signal N_1_2 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO\ : std_logic ;
  signal N_1_3 : std_logic ;
  signal N_1_4 : std_logic ;
  signal N_1_5 : std_logic ;
  signal N_1_6 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349_RETI\ : std_logic ;
  signal N_65771_RETO : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO\ : std_logic ;
  signal N_1_7 : std_logic ;
  signal N_65496_RETI : std_logic ;
  signal N_65775_RETI : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM6_RETI\ : std_logic ;
  signal N_1_8 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_3_RETI\ : std_logic ;
  signal N_1_9 : std_logic ;
  signal N_1_10 : std_logic ;
  signal N_1_11 : std_logic ;
  signal N_1_12 : std_logic ;
  signal N_1_13 : std_logic ;
  signal N_1_14 : std_logic ;
  signal N_1_15 : std_logic ;
  signal N_1_16 : std_logic ;
  signal N_1_17 : std_logic ;
  signal N_1_18 : std_logic ;
  signal N_1_19 : std_logic ;
  signal N_1_20 : std_logic ;
  signal N_1_21 : std_logic ;
  signal N_1_22 : std_logic ;
  signal N_1_23 : std_logic ;
  signal N_1_24 : std_logic ;
  signal N_1_25 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_RETO\ : std_logic ;
  signal N_1_26 : std_logic ;
  signal N_1_27 : std_logic ;
  signal N_1_28 : std_logic ;
  signal N_1_29 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5346_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_0_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7350_RETI\ : std_logic ;
  signal N_1_30 : std_logic ;
  signal N_1_31 : std_logic ;
  signal N_1_32 : std_logic ;
  signal N_1_33 : std_logic ;
  signal N_1_34 : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_I_RETO\ : std_logic ;
  signal N_1_35 : std_logic ;
  signal N_1_36 : std_logic ;
  signal N_1_37 : std_logic ;
  signal N_1_38 : std_logic ;
  signal N_1_39 : std_logic ;
  signal N_1_40 : std_logic ;
  signal N_1_41 : std_logic ;
  signal N_1_42 : std_logic ;
  signal N_1_43 : std_logic ;
  signal N_1_44 : std_logic ;
  signal N_1_45 : std_logic ;
  signal N_1_46 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO\ : std_logic ;
  signal N_1_47 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\ : std_logic ;
  signal N_1_48 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\ : std_logic ;
  signal N_1_49 : std_logic ;
  signal N_1_50 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_TZ_RETO\ : std_logic ;
  signal N_1_51 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO5_RETO\ : std_logic ;
  signal N_1_52 : std_logic ;
  signal N_1_53 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO\ : std_logic ;
  signal N_1_54 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO\ : std_logic ;
  signal N_65609_RETO : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO\ : std_logic ;
  signal N_1_55 : std_logic ;
  signal N_1_56 : std_logic ;
  signal N_59001_RETO : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_RETO\ : std_logic ;
  signal N_58999_RETO : std_logic ;
  signal N_1_57 : std_logic ;
  signal N_59000_RETO : std_logic ;
  signal N_1_58 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_318__G1_RETO\ : std_logic ;
  signal N_1_59 : std_logic ;
  signal RST_RETO : std_logic ;
  signal \GRLFPC2_0.FPO.BUSY_O\ : std_logic ;
  signal N_1_60 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_319__G1_RETO\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_1_RETO\ : std_logic ;
  signal \GRLFPC2_0.FPI.RST_1_RETO\ : std_logic ;
  signal N_1_61 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_372__G1_RETO\ : std_logic ;
  signal N_1_62 : std_logic ;
  signal N_1_63 : std_logic ;
  signal N_2 : std_logic ;
  signal N_3 : std_logic ;
  signal N_4 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\ : std_logic ;
  signal N_65488_RETO : std_logic ;
  signal D_N_7_RETO : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO\ : std_logic ;
  signal N_5 : std_logic ;
  signal N_1_64 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_RETO\ : std_logic ;
  signal N_1_65 : std_logic ;
  signal N_1_66 : std_logic ;
  signal N_1_67 : std_logic ;
  signal N_1_68 : std_logic ;
  signal N_1_69 : std_logic ;
  signal N_1_70 : std_logic ;
  signal N_1_71 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO\ : std_logic ;
  signal N_1_72 : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_RETO\ : std_logic ;
  signal N_1_73 : std_logic ;
  signal N_1_74 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0\ : std_logic ;
  signal \GRLFPC2_0.R.MK.BUSY_RET_0_0_G0_MUX2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4424\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1\ : std_logic ;
  signal N_65609 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7248\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C\ : std_logic ;
  signal N_66444 : std_logic ;
  signal N_66445 : std_logic ;
  signal N_66446 : std_logic ;
  signal N_66563 : std_logic ;
  signal N_66565 : std_logic ;
  signal N_66569 : std_logic ;
  signal N_66571 : std_logic ;
  signal N_66581 : std_logic ;
  signal N_66583 : std_logic ;
  signal N_66585 : std_logic ;
  signal N_66587 : std_logic ;
  signal N_66593 : std_logic ;
  signal N_66595 : std_logic ;
  signal N_66597 : std_logic ;
  signal N_66607 : std_logic ;
  signal N_66615 : std_logic ;
  signal N_66617 : std_logic ;
  signal N_66927 : std_logic ;
  signal N_66928 : std_logic ;
  signal N_66969 : std_logic ;
  signal N_66970 : std_logic ;
  signal N_66971 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_I\ : std_logic ;
  signal N_27258_I : std_logic ;
  signal RST_I : std_logic ;
  signal N_61587_I_0 : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_1_0\ : std_logic ;
  signal \GRLFPC2_0.R.MK.RST2_0\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_0\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_1_1\ : std_logic ;
  signal \GRLFPC2_0.R.MK.RST2_1\ : std_logic ;
  signal \GRLFPC2_0.R.MK.RST_0\ : std_logic ;
  signal \GRLFPC2_0.R.MK.RST_4_0\ : std_logic ;
  signal \GRLFPC2_0.R.MK.RST2_2\ : std_logic ;
  signal \GRLFPC2_0.R.MK.RST2_O_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.ANNULFPU_1_O_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_RETI_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_RETI_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10936_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN13_RESVEC_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10936_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN13_RESVEC_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_3\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_1_2\ : std_logic ;
  signal \GRLFPC2_0.R.MK.RST_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_I_A7_10_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_I_A7_6_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0_N_5_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_1_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0_M3_I_A3_0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0_N_5_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_1_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0_M3_I_A3_0_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM12_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7778_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7777_0\ : std_logic ;
  signal N_65516_0 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM12_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7778_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7777_1\ : std_logic ;
  signal N_65516_1 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\ : std_logic ;
  signal N_65549_0 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN12_SRTOSTICKY_1_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5346_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5346_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_16\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_18\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_19\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_20\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_21\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_22\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_23\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_24\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_16\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_16\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_25\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_26\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_18\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_18\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_27\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_19\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_19\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_28\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_20\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_20\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_29\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_21\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_21\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_30\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_22\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_22\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_31\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_23\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_23\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_32\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_24\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_24\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_33\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_25\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_25\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_34\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_26\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_26\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_35\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_27\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_27\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_36\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_28\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_28\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_37\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_29\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_29\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_38\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_30\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_30\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_39\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_31\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_31\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_40\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_32\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_32\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_41\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_33\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_33\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_42\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_34\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_34\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_43\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_35\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_35\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_44\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_36\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_36\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_45\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_37\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_37\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_46\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_38\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_38\ : std_logic ;
  signal N_65771_RETO_0 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO_0\ : std_logic ;
  signal N_65771_RETO_1 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO_1\ : std_logic ;
  signal N_65771_RETO_2 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO_2\ : std_logic ;
  signal N_65771_RETO_3 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO_3\ : std_logic ;
  signal N_65771_RETO_4 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO_4\ : std_logic ;
  signal N_65771_RETO_5 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO_5\ : std_logic ;
  signal N_65771_RETO_6 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO_6\ : std_logic ;
  signal N_65771_RETO_7 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_2\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_0_0\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_1_1_0\ : std_logic ;
  signal \GRLFPC2_0.R.MK.RST2_1_0\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_0_1\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_1_1_1\ : std_logic ;
  signal \GRLFPC2_0.R.MK.RST2_1_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_2\ : std_logic ;
  signal N_65488_RETO_0 : std_logic ;
  signal N_65488_0 : std_logic ;
  signal D_N_7_RETO_0 : std_logic ;
  signal D_N_7_0 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_0\ : std_logic ;
  signal N_32738_1_0 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10934_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10934_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_513_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_479_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_3\ : std_logic ;
  signal N_65488_1 : std_logic ;
  signal D_N_7_1 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_TZ_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_1_3\ : std_logic ;
  signal \GRLFPC2_0.R.MK.RST2_3\ : std_logic ;
  signal \GRLFPC2_0.V.STATE_2_SQMUXA0\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN1_V.STATE0\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.FSR.FCC80\ : std_logic ;
  signal \GRLFPC2_0.V.FSR.CEXC_2_SQMUXA0\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN1_V.STATE0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_00\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS0\ : std_logic ;
  signal N_6 : std_logic ;
  signal N_7 : std_logic ;
  signal N_8 : std_logic ;
  signal N_9 : std_logic ;
  signal N_10 : std_logic ;
  signal N_11 : std_logic ;
  signal N_12 : std_logic ;
  signal N_13 : std_logic ;
  signal N_14 : std_logic ;
  signal N_15 : std_logic ;
  signal N_16 : std_logic ;
  signal N_17 : std_logic ;
  signal N_18 : std_logic ;
  signal N_19 : std_logic ;
  signal N_20 : std_logic ;
  signal N_21 : std_logic ;
  signal N_22 : std_logic ;
  signal N_23 : std_logic ;
  signal N_24 : std_logic ;
  signal N_25 : std_logic ;
  signal N_26 : std_logic ;
  signal N_27 : std_logic ;
  signal N_28 : std_logic ;
  signal N_29 : std_logic ;
  signal N_30 : std_logic ;
  signal N_31 : std_logic ;
  signal N_32 : std_logic ;
  signal N_33 : std_logic ;
  signal N_34 : std_logic ;
  signal N_35 : std_logic ;
  signal N_36 : std_logic ;
  signal N_37 : std_logic ;
  signal N_38 : std_logic ;
  signal N_39 : std_logic ;
  signal N_40 : std_logic ;
  signal N_41 : std_logic ;
  signal N_42 : std_logic ;
  signal N_43 : std_logic ;
  signal N_44 : std_logic ;
  signal N_45 : std_logic ;
  signal N_46 : std_logic ;
  signal N_47 : std_logic ;
  signal N_48 : std_logic ;
  signal N_49 : std_logic ;
  signal N_50 : std_logic ;
  signal N_51 : std_logic ;
  signal N_52 : std_logic ;
  signal N_53 : std_logic ;
  signal N_54 : std_logic ;
  signal N_55 : std_logic ;
  signal N_56 : std_logic ;
  signal N_57 : std_logic ;
  signal N_58 : std_logic ;
  signal N_59 : std_logic ;
  signal N_60 : std_logic ;
  signal N_61 : std_logic ;
  signal N_62 : std_logic ;
  signal N_63 : std_logic ;
  signal N_64 : std_logic ;
  signal N_65 : std_logic ;
  signal N_66 : std_logic ;
  signal N_67 : std_logic ;
  signal N_68 : std_logic ;
  signal N_69 : std_logic ;
  signal N_70 : std_logic ;
  signal N_71 : std_logic ;
  signal N_72 : std_logic ;
  signal N_73 : std_logic ;
  signal N_74 : std_logic ;
  signal N_75 : std_logic ;
  signal N_76 : std_logic ;
  signal N_77 : std_logic ;
  signal N_78 : std_logic ;
  signal N_79 : std_logic ;
  signal N_80 : std_logic ;
  signal N_81 : std_logic ;
  signal N_82 : std_logic ;
  signal N_83 : std_logic ;
  signal N_84 : std_logic ;
  signal N_85 : std_logic ;
  signal N_86 : std_logic ;
  signal N_87 : std_logic ;
  signal N_88 : std_logic ;
  signal N_89 : std_logic ;
  signal N_90 : std_logic ;
  signal N_91 : std_logic ;
  signal N_92 : std_logic ;
  signal N_93 : std_logic ;
  signal N_94 : std_logic ;
  signal N_95 : std_logic ;
  signal N_96 : std_logic ;
  signal N_97 : std_logic ;
  signal N_98 : std_logic ;
  signal N_99 : std_logic ;
  signal N_100 : std_logic ;
  signal N_101 : std_logic ;
  signal N_102 : std_logic ;
  signal N_103 : std_logic ;
  signal N_104 : std_logic ;
  signal N_105 : std_logic ;
  signal N_106 : std_logic ;
  signal N_107 : std_logic ;
  signal N_108 : std_logic ;
  signal N_109 : std_logic ;
  signal N_110 : std_logic ;
  signal N_111 : std_logic ;
  signal N_112 : std_logic ;
  signal N_113 : std_logic ;
  signal N_114 : std_logic ;
  signal N_115 : std_logic ;
  signal N_116 : std_logic ;
  signal N_117 : std_logic ;
  signal N_118 : std_logic ;
  signal N_119 : std_logic ;
  signal N_120 : std_logic ;
  signal N_121 : std_logic ;
  signal N_122 : std_logic ;
  signal N_123 : std_logic ;
  signal N_124 : std_logic ;
  signal N_125 : std_logic ;
  signal N_126 : std_logic ;
  signal N_127 : std_logic ;
  signal N_128 : std_logic ;
  signal N_129 : std_logic ;
  signal N_130 : std_logic ;
  signal N_131 : std_logic ;
  signal N_132 : std_logic ;
  signal N_133 : std_logic ;
  signal N_134 : std_logic ;
  signal N_135 : std_logic ;
  signal N_136 : std_logic ;
  signal N_137 : std_logic ;
  signal N_138 : std_logic ;
  signal N_139 : std_logic ;
  signal N_140 : std_logic ;
  signal N_141 : std_logic ;
  signal N_142 : std_logic ;
  signal N_143 : std_logic ;
  signal N_144 : std_logic ;
  signal N_145 : std_logic ;
  signal N_146 : std_logic ;
  signal N_147 : std_logic ;
  signal N_148 : std_logic ;
  signal N_149 : std_logic ;
  signal N_150 : std_logic ;
  signal N_151 : std_logic ;
  signal N_152 : std_logic ;
  signal N_153 : std_logic ;
  signal N_154 : std_logic ;
  signal N_155 : std_logic ;
  signal N_156 : std_logic ;
  signal N_157 : std_logic ;
  signal N_158 : std_logic ;
  signal N_159 : std_logic ;
  signal N_160 : std_logic ;
  signal N_161 : std_logic ;
  signal N_162 : std_logic ;
  signal N_163 : std_logic ;
  signal N_164 : std_logic ;
  signal N_165 : std_logic ;
  signal N_166 : std_logic ;
  signal N_167 : std_logic ;
  signal N_168 : std_logic ;
  signal N_169 : std_logic ;
  signal N_170 : std_logic ;
  signal N_171 : std_logic ;
  signal N_172 : std_logic ;
  signal N_173 : std_logic ;
  signal N_174 : std_logic ;
  signal N_175 : std_logic ;
  signal N_176 : std_logic ;
  signal N_177 : std_logic ;
  signal N_178 : std_logic ;
  signal N_179 : std_logic ;
  signal N_180 : std_logic ;
  signal N_181 : std_logic ;
  signal N_182 : std_logic ;
  signal N_183 : std_logic ;
  signal N_184 : std_logic ;
  signal N_185 : std_logic ;
  signal N_186 : std_logic ;
  signal N_187 : std_logic ;
  signal N_188 : std_logic ;
  signal N_189 : std_logic ;
  signal N_190 : std_logic ;
  signal N_191 : std_logic ;
  signal N_192 : std_logic ;
  signal N_193 : std_logic ;
  signal N_194 : std_logic ;
  signal N_195 : std_logic ;
  signal N_196 : std_logic ;
  signal N_197 : std_logic ;
  signal N_198 : std_logic ;
  signal N_199 : std_logic ;
  signal N_200 : std_logic ;
  signal N_201 : std_logic ;
  signal N_202 : std_logic ;
  signal N_203 : std_logic ;
  signal N_204 : std_logic ;
  signal N_205 : std_logic ;
  signal N_206 : std_logic ;
  signal N_207 : std_logic ;
  signal N_208 : std_logic ;
  signal N_209 : std_logic ;
  signal N_210 : std_logic ;
  signal N_211 : std_logic ;
  signal N_212 : std_logic ;
  signal N_213 : std_logic ;
  signal N_214 : std_logic ;
  signal N_215 : std_logic ;
  signal N_216 : std_logic ;
  signal N_217 : std_logic ;
  signal N_218 : std_logic ;
  signal N_219 : std_logic ;
  signal N_220 : std_logic ;
  signal N_221 : std_logic ;
  signal N_222 : std_logic ;
  signal N_223 : std_logic ;
  signal N_224 : std_logic ;
  signal N_225 : std_logic ;
  signal N_226 : std_logic ;
  signal N_227 : std_logic ;
  signal N_228 : std_logic ;
  signal N_229 : std_logic ;
  signal N_230 : std_logic ;
  signal N_231 : std_logic ;
  signal N_232 : std_logic ;
  signal N_233 : std_logic ;
  signal N_234 : std_logic ;
  signal N_235 : std_logic ;
  signal N_236 : std_logic ;
  signal N_237 : std_logic ;
  signal N_238 : std_logic ;
  signal N_239 : std_logic ;
  signal N_240 : std_logic ;
  signal N_241 : std_logic ;
  signal N_242 : std_logic ;
  signal N_243 : std_logic ;
  signal N_244 : std_logic ;
  signal N_245 : std_logic ;
  signal N_246 : std_logic ;
  signal N_247 : std_logic ;
  signal N_248 : std_logic ;
  signal N_249 : std_logic ;
  signal N_250 : std_logic ;
  signal N_251 : std_logic ;
  signal N_252 : std_logic ;
  signal N_253 : std_logic ;
  signal N_254 : std_logic ;
  signal N_255 : std_logic ;
  signal N_256 : std_logic ;
  signal N_257 : std_logic ;
  signal N_258 : std_logic ;
  signal N_259 : std_logic ;
  signal N_260 : std_logic ;
  signal N_261 : std_logic ;
  signal N_262 : std_logic ;
  signal N_263 : std_logic ;
  signal N_264 : std_logic ;
  signal N_265 : std_logic ;
  signal N_266 : std_logic ;
  signal N_267 : std_logic ;
  signal N_268 : std_logic ;
  signal N_269 : std_logic ;
  signal N_270 : std_logic ;
  signal N_271 : std_logic ;
  signal N_272 : std_logic ;
  signal N_273 : std_logic ;
  signal N_274 : std_logic ;
  signal N_275 : std_logic ;
  signal N_276 : std_logic ;
  signal N_277 : std_logic ;
  signal N_278 : std_logic ;
  signal N_279 : std_logic ;
  signal N_280 : std_logic ;
  signal N_281 : std_logic ;
  signal N_282 : std_logic ;
  signal N_283 : std_logic ;
  signal N_284 : std_logic ;
  signal N_285 : std_logic ;
  signal N_286 : std_logic ;
  signal N_287 : std_logic ;
  signal N_288 : std_logic ;
  signal N_289 : std_logic ;
  signal N_290 : std_logic ;
  signal N_291 : std_logic ;
  signal N_292 : std_logic ;
  signal N_293 : std_logic ;
  signal N_294 : std_logic ;
  signal N_295 : std_logic ;
  signal N_296 : std_logic ;
  signal N_297 : std_logic ;
  signal N_298 : std_logic ;
  signal N_299 : std_logic ;
  signal N_300 : std_logic ;
  signal N_301 : std_logic ;
  signal N_302 : std_logic ;
  signal N_303 : std_logic ;
  signal N_304 : std_logic ;
  signal N_305 : std_logic ;
  signal N_306 : std_logic ;
  signal N_307 : std_logic ;
  signal N_308 : std_logic ;
  signal N_309 : std_logic ;
  signal N_310 : std_logic ;
  signal N_311 : std_logic ;
  signal N_312 : std_logic ;
  signal N_313 : std_logic ;
  signal N_314 : std_logic ;
  signal N_315 : std_logic ;
  signal N_316 : std_logic ;
  signal N_317 : std_logic ;
  signal N_318 : std_logic ;
  signal N_319 : std_logic ;
  signal N_320 : std_logic ;
  signal N_321 : std_logic ;
  signal N_322 : std_logic ;
  signal N_323 : std_logic ;
  signal N_324 : std_logic ;
  signal N_325 : std_logic ;
  signal N_326 : std_logic ;
  signal N_327 : std_logic ;
  signal N_328 : std_logic ;
  signal N_329 : std_logic ;
  signal N_330 : std_logic ;
  signal N_331 : std_logic ;
  signal N_332 : std_logic ;
  signal N_333 : std_logic ;
  signal N_334 : std_logic ;
  signal N_335 : std_logic ;
  signal N_336 : std_logic ;
  signal N_337 : std_logic ;
  signal N_338 : std_logic ;
  signal N_339 : std_logic ;
  signal N_340 : std_logic ;
  signal N_341 : std_logic ;
  signal N_342 : std_logic ;
  signal N_343 : std_logic ;
  signal N_344 : std_logic ;
  signal N_345 : std_logic ;
  signal N_346 : std_logic ;
  signal N_347 : std_logic ;
  signal N_348 : std_logic ;
  signal N_349 : std_logic ;
  signal N_350 : std_logic ;
  signal N_351 : std_logic ;
  signal N_352 : std_logic ;
  signal N_353 : std_logic ;
  signal N_354 : std_logic ;
  signal N_355 : std_logic ;
  signal N_356 : std_logic ;
  signal N_357 : std_logic ;
  signal N_358 : std_logic ;
  signal N_359 : std_logic ;
  signal N_360 : std_logic ;
  signal N_361 : std_logic ;
  signal N_362 : std_logic ;
  signal N_363 : std_logic ;
  signal N_364 : std_logic ;
  signal N_365 : std_logic ;
  signal N_366 : std_logic ;
  signal N_367 : std_logic ;
  signal N_368 : std_logic ;
  signal N_369 : std_logic ;
  signal N_370 : std_logic ;
  signal N_371 : std_logic ;
  signal N_372 : std_logic ;
  signal N_373 : std_logic ;
  signal N_374 : std_logic ;
  signal N_375 : std_logic ;
  signal N_376 : std_logic ;
  signal N_377 : std_logic ;
  signal N_378 : std_logic ;
  signal N_379 : std_logic ;
  signal N_380 : std_logic ;
  signal N_381 : std_logic ;
  signal N_382 : std_logic ;
  signal N_383 : std_logic ;
  signal N_384 : std_logic ;
  signal N_385 : std_logic ;
  signal N_386 : std_logic ;
  signal N_387 : std_logic ;
  signal N_388 : std_logic ;
  signal N_389 : std_logic ;
  signal N_390 : std_logic ;
  signal N_391 : std_logic ;
  signal N_392 : std_logic ;
  signal N_393 : std_logic ;
  signal N_394 : std_logic ;
  signal N_395 : std_logic ;
  signal N_396 : std_logic ;
  signal N_397 : std_logic ;
  signal N_398 : std_logic ;
  signal N_399 : std_logic ;
  signal N_400 : std_logic ;
  signal N_401 : std_logic ;
  signal N_402 : std_logic ;
  signal N_403 : std_logic ;
  signal N_404 : std_logic ;
  signal N_405 : std_logic ;
  signal N_406 : std_logic ;
  signal N_407 : std_logic ;
  signal N_408 : std_logic ;
  signal N_409 : std_logic ;
  signal N_410 : std_logic ;
  signal N_411 : std_logic ;
  signal N_412 : std_logic ;
  signal N_413 : std_logic ;
  signal N_414 : std_logic ;
  signal N_415 : std_logic ;
  signal N_416 : std_logic ;
  signal N_417 : std_logic ;
  signal N_418 : std_logic ;
  signal N_419 : std_logic ;
  signal N_420 : std_logic ;
  signal N_421 : std_logic ;
  signal N_422 : std_logic ;
  signal N_423 : std_logic ;
  signal N_424 : std_logic ;
  signal N_425 : std_logic ;
  signal N_426 : std_logic ;
  signal N_427 : std_logic ;
  signal N_428 : std_logic ;
  signal N_429 : std_logic ;
  signal N_430 : std_logic ;
  signal N_431 : std_logic ;
  signal N_432 : std_logic ;
  signal N_433 : std_logic ;
  signal N_434 : std_logic ;
  signal N_435 : std_logic ;
  signal N_436 : std_logic ;
  signal N_437 : std_logic ;
  signal N_0 : std_logic ;
  signal N_1_75 : std_logic ;
  signal N_2_0 : std_logic ;
  signal N_3_0 : std_logic ;
  signal N_4_0 : std_logic ;
  signal N_5_0 : std_logic ;
  signal N_6_0 : std_logic ;
  signal N_7_0 : std_logic ;
  signal N_8_0 : std_logic ;
  signal N_9_0 : std_logic ;
  signal N_10_0 : std_logic ;
  signal N_11_0 : std_logic ;
  signal N_12_0 : std_logic ;
  signal N_13_0 : std_logic ;
  signal N_14_0 : std_logic ;
  signal N_15_0 : std_logic ;
  signal N_16_0 : std_logic ;
  signal N_17_0 : std_logic ;
  signal N_18_0 : std_logic ;
  signal N_19_0 : std_logic ;
  signal N_20_0 : std_logic ;
  signal N_21_0 : std_logic ;
  signal N_22_0 : std_logic ;
  signal N_23_0 : std_logic ;
  signal N_24_0 : std_logic ;
  signal N_25_0 : std_logic ;
  signal N_26_0 : std_logic ;
  signal N_27_0 : std_logic ;
  signal N_28_0 : std_logic ;
  signal N_29_0 : std_logic ;
  signal N_30_0 : std_logic ;
  signal N_31_0 : std_logic ;
  signal N_32_0 : std_logic ;
  signal N_33_0 : std_logic ;
  signal N_34_0 : std_logic ;
  signal N_35_0 : std_logic ;
  signal N_36_0 : std_logic ;
  signal N_37_0 : std_logic ;
  signal N_38_0 : std_logic ;
  signal N_39_0 : std_logic ;
  signal N_40_0 : std_logic ;
  signal N_41_0 : std_logic ;
  signal N_42_0 : std_logic ;
  signal N_43_0 : std_logic ;
  signal N_44_0 : std_logic ;
  signal N_45_0 : std_logic ;
  signal N_46_0 : std_logic ;
  signal N_47_0 : std_logic ;
  signal N_48_0 : std_logic ;
  signal N_49_0 : std_logic ;
  signal N_50_0 : std_logic ;
  signal N_51_0 : std_logic ;
  signal N_52_0 : std_logic ;
  signal N_53_0 : std_logic ;
  signal N_54_0 : std_logic ;
  signal N_55_0 : std_logic ;
  signal N_56_0 : std_logic ;
  signal N_57_0 : std_logic ;
  signal N_58_0 : std_logic ;
  signal N_59_0 : std_logic ;
  signal N_60_0 : std_logic ;
  signal N_61_0 : std_logic ;
  signal N_62_0 : std_logic ;
  signal N_63_0 : std_logic ;
  signal N_64_0 : std_logic ;
  signal N_65_0 : std_logic ;
  signal N_66_0 : std_logic ;
  signal N_67_0 : std_logic ;
  signal N_68_0 : std_logic ;
  signal N_69_0 : std_logic ;
  signal N_70_0 : std_logic ;
  signal N_71_0 : std_logic ;
  signal N_72_0 : std_logic ;
  signal N_73_0 : std_logic ;
  signal N_74_0 : std_logic ;
  signal N_75_0 : std_logic ;
  signal N_76_0 : std_logic ;
  signal N_77_0 : std_logic ;
  signal N_78_0 : std_logic ;
  signal N_79_0 : std_logic ;
  signal N_80_0 : std_logic ;
  signal N_81_0 : std_logic ;
  signal N_82_0 : std_logic ;
  signal N_83_0 : std_logic ;
  signal N_84_0 : std_logic ;
  signal N_85_0 : std_logic ;
  signal N_86_0 : std_logic ;
  signal N_87_0 : std_logic ;
  signal N_88_0 : std_logic ;
  signal N_89_0 : std_logic ;
  signal N_90_0 : std_logic ;
  signal N_91_0 : std_logic ;
  signal N_92_0 : std_logic ;
  signal N_93_0 : std_logic ;
  signal N_94_0 : std_logic ;
  signal N_95_0 : std_logic ;
  signal N_96_0 : std_logic ;
  signal N_97_0 : std_logic ;
  signal N_98_0 : std_logic ;
  signal N_99_0 : std_logic ;
  signal N_100_0 : std_logic ;
  signal N_101_0 : std_logic ;
  signal N_102_0 : std_logic ;
  signal N_103_0 : std_logic ;
  signal N_104_0 : std_logic ;
  signal N_105_0 : std_logic ;
  signal N_106_0 : std_logic ;
  signal N_107_0 : std_logic ;
  signal N_108_0 : std_logic ;
  signal N_109_0 : std_logic ;
  signal N_110_0 : std_logic ;
  signal N_111_0 : std_logic ;
  signal N_112_0 : std_logic ;
  signal N_113_0 : std_logic ;
  signal N_114_0 : std_logic ;
  signal N_115_0 : std_logic ;
  signal N_116_0 : std_logic ;
  signal N_117_0 : std_logic ;
  signal N_118_0 : std_logic ;
  signal N_119_0 : std_logic ;
  signal N_120_0 : std_logic ;
  signal N_121_0 : std_logic ;
  signal N_122_0 : std_logic ;
  signal N_123_0 : std_logic ;
  signal N_124_0 : std_logic ;
  signal N_125_0 : std_logic ;
  signal N_126_0 : std_logic ;
  signal N_127_0 : std_logic ;
  signal N_128_0 : std_logic ;
  signal N_129_0 : std_logic ;
  signal N_130_0 : std_logic ;
  signal N_131_0 : std_logic ;
  signal N_132_0 : std_logic ;
  signal N_133_0 : std_logic ;
  signal N_134_0 : std_logic ;
  signal N_135_0 : std_logic ;
  signal N_136_0 : std_logic ;
  signal N_137_0 : std_logic ;
  signal N_138_0 : std_logic ;
  signal N_139_0 : std_logic ;
  signal N_140_0 : std_logic ;
  signal N_141_0 : std_logic ;
  signal N_142_0 : std_logic ;
  signal N_143_0 : std_logic ;
  signal N_144_0 : std_logic ;
  signal N_145_0 : std_logic ;
  signal N_146_0 : std_logic ;
  signal N_147_0 : std_logic ;
  signal N_148_0 : std_logic ;
  signal N_149_0 : std_logic ;
  signal N_150_0 : std_logic ;
  signal N_151_0 : std_logic ;
  signal N_152_0 : std_logic ;
  signal N_153_0 : std_logic ;
  signal N_154_0 : std_logic ;
  signal N_155_0 : std_logic ;
  signal N_156_0 : std_logic ;
  signal N_157_0 : std_logic ;
  signal N_158_0 : std_logic ;
  signal N_159_0 : std_logic ;
  signal N_160_0 : std_logic ;
  signal N_161_0 : std_logic ;
  signal N_162_0 : std_logic ;
  signal N_163_0 : std_logic ;
  signal N_602 : std_logic ;
  signal N_603 : std_logic ;
  signal N_604 : std_logic ;
  signal N_605 : std_logic ;
  signal N_606 : std_logic ;
  signal N_607 : std_logic ;
  signal N_608 : std_logic ;
  signal N_609 : std_logic ;
  signal N_610 : std_logic ;
  signal N_611 : std_logic ;
  signal N_612 : std_logic ;
  signal N_613 : std_logic ;
  signal N_614 : std_logic ;
  signal N_615 : std_logic ;
  signal N_616 : std_logic ;
  signal N_617 : std_logic ;
  signal N_618 : std_logic ;
  signal N_619 : std_logic ;
  signal N_620 : std_logic ;
  signal N_621 : std_logic ;
  signal N_622 : std_logic ;
  signal N_623 : std_logic ;
  signal N_624 : std_logic ;
  signal N_625 : std_logic ;
  signal N_626 : std_logic ;
  signal N_627 : std_logic ;
  signal N_628 : std_logic ;
  signal N_629 : std_logic ;
  signal N_630 : std_logic ;
  signal N_631 : std_logic ;
  signal N_632 : std_logic ;
  signal N_633 : std_logic ;
  signal N_634 : std_logic ;
  signal N_635 : std_logic ;
  signal N_636 : std_logic ;
  signal N_637 : std_logic ;
  signal N_638 : std_logic ;
  signal N_639 : std_logic ;
  signal N_640 : std_logic ;
  signal N_641 : std_logic ;
  signal N_642 : std_logic ;
  signal N_643 : std_logic ;
  signal N_644 : std_logic ;
  signal N_645 : std_logic ;
  signal N_646 : std_logic ;
  signal N_647 : std_logic ;
  signal N_648 : std_logic ;
  signal N_649 : std_logic ;
  signal N_650 : std_logic ;
  signal N_651 : std_logic ;
  signal N_652 : std_logic ;
  signal N_653 : std_logic ;
  signal N_654 : std_logic ;
  signal N_655 : std_logic ;
  signal N_656 : std_logic ;
  signal N_657 : std_logic ;
  signal N_658 : std_logic ;
  signal N_659 : std_logic ;
  signal N_660 : std_logic ;
  signal N_661 : std_logic ;
  signal N_662 : std_logic ;
  signal N_663 : std_logic ;
  signal N_664 : std_logic ;
  signal N_665 : std_logic ;
  signal N_666 : std_logic ;
  signal N_667 : std_logic ;
  signal N_668 : std_logic ;
  signal N_669 : std_logic ;
  signal N_670 : std_logic ;
  signal N_671 : std_logic ;
  signal N_672 : std_logic ;
  signal N_673 : std_logic ;
  signal N_674 : std_logic ;
  signal N_675 : std_logic ;
  signal N_676 : std_logic ;
  signal N_677 : std_logic ;
  signal N_678 : std_logic ;
  signal N_679 : std_logic ;
  signal N_680 : std_logic ;
  signal N_681 : std_logic ;
  signal N_682 : std_logic ;
  signal N_683 : std_logic ;
  signal N_684 : std_logic ;
  signal N_685 : std_logic ;
  signal N_686 : std_logic ;
  signal N_687 : std_logic ;
  signal N_688 : std_logic ;
  signal N_689 : std_logic ;
  signal N_690 : std_logic ;
  signal N_691 : std_logic ;
  signal N_692 : std_logic ;
  signal N_693 : std_logic ;
  signal N_694 : std_logic ;
  signal N_695 : std_logic ;
  signal N_696 : std_logic ;
  signal N_697 : std_logic ;
  signal N_698 : std_logic ;
  signal N_699 : std_logic ;
  signal N_700 : std_logic ;
  signal N_701 : std_logic ;
  signal N_702 : std_logic ;
  signal N_703 : std_logic ;
  signal N_704 : std_logic ;
  signal N_705 : std_logic ;
  signal N_706 : std_logic ;
  signal N_707 : std_logic ;
  signal N_708 : std_logic ;
  signal N_709 : std_logic ;
  signal N_710 : std_logic ;
  signal N_711 : std_logic ;
  signal N_712 : std_logic ;
  signal N_713 : std_logic ;
  signal N_714 : std_logic ;
  signal N_715 : std_logic ;
  signal N_716 : std_logic ;
  signal N_717 : std_logic ;
  signal N_718 : std_logic ;
  signal N_719 : std_logic ;
  signal N_720 : std_logic ;
  signal N_721 : std_logic ;
  signal N_722 : std_logic ;
  signal N_723 : std_logic ;
  signal N_724 : std_logic ;
  signal N_725 : std_logic ;
  signal N_726 : std_logic ;
  signal N_727 : std_logic ;
  signal N_728 : std_logic ;
  signal N_729 : std_logic ;
  signal CPO_EXCZ : std_logic ;
  signal CPO_CCVZ : std_logic ;
  signal CPO_LDLOCKZ : std_logic ;
  signal CPO_HOLDNZ : std_logic ;
  signal RFI1_REN1Z : std_logic ;
  signal RFI1_REN2Z : std_logic ;
  signal RFI1_WRENZ : std_logic ;
  signal RFI2_REN1Z : std_logic ;
  signal RFI2_REN2Z : std_logic ;
  signal RFI2_WRENZ : std_logic ;
begin
VCC <= '1';
GND <= '0';
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIFMH6_0_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"000000aa0000aa55")
port map (
sumout => N_27260,
cout => N_29683,
shareout => N_29684,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(29),
cin => GND,
sharein => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIMI0Q_30_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000fcc00000c33c")
port map (
sumout => N_27262,
cout => N_29686,
shareout => N_29687,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(29),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(30),
cin => N_29683,
sharein => N_29684);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIGHES1_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27264,
cout => N_29689,
shareout => N_29690,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(31),
cin => N_29686,
sharein => N_29687);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI6FA14_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27266,
cout => N_29692,
shareout => N_29693,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(32),
cin => N_29689,
sharein => N_29690);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIKA2B8_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27268,
cout => N_29695,
shareout => N_29696,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(33),
cin => N_29692,
sharein => N_29693);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNII1IUG_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27270,
cout => N_29698,
shareout => N_29699,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(34),
cin => N_29695,
sharein => N_29696);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIGFH521_35_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27272,
cout => N_29701,
shareout => N_29702,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(35),
cin => N_29698,
sharein => N_29699);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIEBGJ42_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27274,
cout => N_29704,
shareout => N_29705,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(36),
cin => N_29701,
sharein => N_29702);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIC3EF94_37_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27276,
cout => N_29707,
shareout => N_29708,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(37),
cin => N_29704,
sharein => N_29705);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIAJ97J8_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27278,
cout => N_29710,
shareout => N_29711,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(38),
cin => N_29707,
sharein => N_29708);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI8J0N6H_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27280,
cout => N_29713,
shareout => N_29714,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(39),
cin => N_29710,
sharein => N_29711);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIOQEMD21_40_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27282,
cout => N_29716,
shareout => N_29717,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(40),
cin => N_29713,
sharein => N_29714);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIQ9BLR42_41_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27284,
cout => N_29719,
shareout => N_29720,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(41),
cin => N_29716,
sharein => N_29717);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI084JN9_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27286,
cout => N_29722,
shareout => N_29723,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(42),
cin => N_29719,
sharein => N_29720);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIE4MEFJ_43_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27288,
cout => N_29725,
shareout => N_29726,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(43),
cin => N_29722,
sharein => N_29723);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNICTP5V61_44_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27290,
cout => N_29728,
shareout => N_29729,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(44),
cin => N_29725,
sharein => N_29726);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNINGLD0E2_45_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27292,
cout => N_29731,
shareout => N_29732,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(45),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(45),
cin => N_29728,
sharein => N_29729);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI2MO31S_46_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27294,
cout => N_29734,
shareout => N_29735,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(46),
cin => N_29731,
sharein => N_29732);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIQ0VF2O1_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27296,
cout => N_29737,
shareout => N_29738,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(47),
cin => N_29734,
sharein => N_29735);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNICMB85G3_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27298,
cout => N_29740,
shareout => N_29741,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(48),
cin => N_29737,
sharein => N_29738);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNII15PA03_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27300,
cout => N_29743,
shareout => N_29744,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(49),
cin => N_29740,
sharein => N_29741);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIIVNQL02_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27302,
cout => N_29746,
shareout => N_29747,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(50),
cin => N_29743,
sharein => N_29744);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIKRTTB1_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27304,
cout => N_29749,
shareout => N_29750,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(51),
cin => N_29746,
sharein => N_29747);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIQJ94O2_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27306,
cout => N_29752,
shareout => N_29753,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(52),
cin => N_29749,
sharein => N_29750);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI841HG5_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27308,
cout => N_29755,
shareout => N_29756,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(53),
cin => N_29752,
sharein => N_29753);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI65GA1B_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27310,
cout => N_29758,
shareout => N_29759,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(54),
cin => N_29755,
sharein => N_29756);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI47ET2M_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27312,
cout => N_29761,
shareout => N_29762,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(55),
cin => N_29758,
sharein => N_29759);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI2BA36C1_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27314,
cout => N_29764,
shareout => N_29765,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(56),
cin => N_29761,
sharein => N_29762);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI0J2FCO2_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27316,
cout => N_6,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(57),
cin => N_29764,
sharein => N_29765);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIFMH6_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27259,
cout => N_29770,
shareout => N_29771,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(29),
cin => GND,
sharein => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI0PGL_30_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27261,
cout => N_29773,
shareout => N_29774,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(30),
cin => N_29770,
sharein => N_29771);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI4UEJ1_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27263,
cout => N_29776,
shareout => N_29777,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(31),
cin => N_29773,
sharein => N_29774);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIE8BF3_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27265,
cout => N_29779,
shareout => N_29780,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(32),
cin => N_29776,
sharein => N_29777);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI4T377_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27267,
cout => N_29782,
shareout => N_29783,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(33),
cin => N_29779,
sharein => N_29780);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNII6LME_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27269,
cout => N_29785,
shareout => N_29786,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(34),
cin => N_29782,
sharein => N_29783);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIGPNLT_35_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27271,
cout => N_29788,
shareout => N_29789,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(35),
cin => N_29785,
sharein => N_29786);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIEVSJR1_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27273,
cout => N_29791,
shareout => N_29792,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(36),
cin => N_29788,
sharein => N_29789);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNICB7GN3_37_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27275,
cout => N_29794,
shareout => N_29795,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(37),
cin => N_29791,
sharein => N_29792);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIA3S8F7_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27277,
cout => N_29797,
shareout => N_29798,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(38),
cin => N_29794,
sharein => N_29795);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI8J5QUE_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27279,
cout => N_29800,
shareout => N_29801,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(39),
cin => N_29797,
sharein => N_29798);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIOQOSTT_40_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27281,
cout => N_29803,
shareout => N_29804,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(40),
cin => N_29800,
sharein => N_29801);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIQ9V1SR1_41_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27283,
cout => N_29806,
shareout => N_29807,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(41),
cin => N_29803,
sharein => N_29804);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI08CCON3_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27285,
cout => N_29809,
shareout => N_29810,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(42),
cin => N_29806,
sharein => N_29807);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIE461HF3_43_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27287,
cout => N_29812,
shareout => N_29813,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(43),
cin => N_29809,
sharein => N_29810);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNICTPA2V2_44_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27289,
cout => N_29815,
shareout => N_29816,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(44),
cin => N_29812,
sharein => N_29813);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNINGLN6U1_45_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27291,
cout => N_29818,
shareout => N_29819,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(45),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(45),
cin => N_29815,
sharein => N_29816);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI2MONDS3_46_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27293,
cout => N_29821,
shareout => N_29822,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(46),
cin => N_29818,
sharein => N_29819);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIQ0VNRO3_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27295,
cout => N_29824,
shareout => N_29825,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(47),
cin => N_29821,
sharein => N_29822);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNICMBONH3_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27297,
cout => N_29827,
shareout => N_29828,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(48),
cin => N_29824,
sharein => N_29825);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNII15PF33_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27299,
cout => N_29830,
shareout => N_29831,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(49),
cin => N_29827,
sharein => N_29828);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIIVNQV62_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27301,
cout => N_29833,
shareout => N_29834,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(50),
cin => N_29830,
sharein => N_29831);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIKRTTVD_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27303,
cout => N_29836,
shareout => N_29837,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(51),
cin => N_29833,
sharein => N_29834);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIQJ940S_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27305,
cout => N_29839,
shareout => N_29840,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(52),
cin => N_29836,
sharein => N_29837);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI841H0O1_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27307,
cout => N_29842,
shareout => N_29843,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(53),
cin => N_29839,
sharein => N_29840);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI65GA1G3_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27309,
cout => N_29845,
shareout => N_29846,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(54),
cin => N_29842,
sharein => N_29843);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI47ET203_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27311,
cout => N_29848,
shareout => N_29849,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(55),
cin => N_29845,
sharein => N_29846);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI2BA3602_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => N_27313,
cout => N_29851,
shareout => N_29852,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(56),
cin => N_29848,
sharein => N_29849);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI0J2FC_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => N_27315,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(57),
cin => N_29851,
sharein => N_29852);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIGOS52_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000ee8800009966")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(0),
cout => N_29857,
shareout => N_29858,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5410\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10552\,
cin => GND,
sharein => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI3BEM5_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(1),
cout => N_29860,
shareout => N_29861,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5391\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(1),
cin => N_29857,
sharein => N_29858);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIUM09D_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(2),
cout => N_29863,
shareout => N_29864,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(2),
cin => N_29860,
sharein => N_29861);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNICLINQ_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(3),
cout => N_29866,
shareout => N_29867,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(3),
cin => N_29863,
sharein => N_29864);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIC39BN1_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(4),
cout => N_29869,
shareout => N_29870,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(4),
cin => N_29866,
sharein => N_29867);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNICU3SE3_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(5),
cout => N_29872,
shareout => N_29873,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(5),
cin => N_29869,
sharein => N_29870);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIESPTT6_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(6),
cout => N_29875,
shareout => N_29876,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(6),
cin => N_29872,
sharein => N_29873);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIK061SD_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(7),
cout => N_29878,
shareout => N_29879,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(7),
cin => N_29875,
sharein => N_29876);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI2HU7OR_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(8),
cout => N_29881,
shareout => N_29882,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(8),
cin => N_29878,
sharein => N_29879);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI0QFLGN1_9_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(9),
cout => N_29884,
shareout => N_29885,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(9),
cin => N_29881,
sharein => N_29882);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIMFCJ1F3_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(10),
cout => N_29887,
shareout => N_29888,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(10),
cin => N_29884,
sharein => N_29885);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI4R5F3U2_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(11),
cout => N_29890,
shareout => N_29891,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(11),
cin => N_29887,
sharein => N_29888);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI2IO67S1_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(12),
cout => N_29893,
shareout => N_29894,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(12),
cin => N_29890,
sharein => N_29891);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI00ULEO3_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(13),
cout => N_29896,
shareout => N_29897,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(13),
cin => N_29893,
sharein => N_29894);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIUR8KTG3_14_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(14),
cout => N_29899,
shareout => N_29900,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(14),
cin => N_29896,
sharein => N_29897);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNISJUGR13_15_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(15),
cout => N_29902,
shareout => N_29903,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(15),
cin => N_29899,
sharein => N_29900);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIQ3AAN32_16_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(16),
cout => N_29905,
shareout => N_29906,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(16),
cin => N_29902,
sharein => N_29903);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIO31TE7_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(17),
cout => N_29908,
shareout => N_29909,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(17),
cin => N_29905,
sharein => N_29906);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIM3F2UE_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(18),
cout => N_29911,
shareout => N_29912,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(18),
cin => N_29908,
sharein => N_29909);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIK3BDST_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(19),
cout => N_29914,
shareout => N_29915,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(19),
cin => N_29911,
sharein => N_29912);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI4B33PR1_20_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(20),
cout => N_29917,
shareout => N_29918,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(20),
cin => N_29914,
sharein => N_29915);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI6QJEIN3_21_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(21),
cout => N_29920,
shareout => N_29921,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(21),
cin => N_29917,
sharein => N_29918);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNICOK55F3_22_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(22),
cout => N_29923,
shareout => N_29924,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(22),
cin => N_29920,
sharein => N_29921);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIQKMJAU2_23_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(23),
cout => N_29926,
shareout => N_29927,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(23),
cin => N_29923,
sharein => N_29924);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIODQFLS1_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(24),
cout => N_29929,
shareout => N_29930,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(24),
cin => N_29926,
sharein => N_29927);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIMV18BP3_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(25),
cout => N_29932,
shareout => N_29933,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(25),
cin => N_29929,
sharein => N_29930);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIK3HOMI3_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(26),
cout => N_29935,
shareout => N_29936,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(26),
cin => N_29932,
sharein => N_29933);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIIBFPD53_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000f00000000ff0")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(27),
cout => N_29938,
shareout => N_29939,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(27),
cin => N_29935,
sharein => N_29936);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIGRBRRA2_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000aa00000055aa")
port map (
sumout => \GRLFPC2_0.FPO.FRAC\(28),
cout => N_29941,
shareout => N_29942,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(28),
cin => N_29938,
sharein => N_29939);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI0NNMNL_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "on",
    extended_lut => "off",
    lut_mask => X"0000000000000000")
port map (
sumout => N_27258,
cout => N_7,
cin => N_29941,
sharein => N_29942);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_9_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_10\(47),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9.Z_CARRY_0\,
dataf => N_52273,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(321),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52267);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_9_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_67\(46),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9.Z_CARRY_1\,
dataf => N_52279,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_9\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_9_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_124\(45),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9.Z_CARRY_2\,
dataf => N_52280,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_66\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_9_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(9),
cout => N_52265,
dataf => N_52288,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_123\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_8_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_9\(48),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8.Z_CARRY_0\,
dataf => N_52296,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(320),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52263);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_8_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_66\(47),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8.Z_CARRY_1\,
dataf => N_52302,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_8\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_8_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_123\(46),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8.Z_CARRY_2\,
dataf => N_52303,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_65\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_8_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(8),
cout => N_52261,
dataf => N_52311,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_122\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_24_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_25\(32),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24.Z_CARRY_0\,
dataf => N_52319,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(336),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52259);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_24_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_82\(31),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24.Z_CARRY_1\,
dataf => N_52325,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_24\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_24_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_139\(30),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24.Z_CARRY_2\,
dataf => N_52326,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_81\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_24_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(24),
cout => N_52257,
dataf => N_52334,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_138\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_23_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_24\(33),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23.Z_CARRY_0\,
dataf => N_52342,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(335),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52255);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_23_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_81\(32),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23.Z_CARRY_1\,
dataf => N_52348,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_23\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_23_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_138\(31),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23.Z_CARRY_2\,
dataf => N_52349,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_80\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_23_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(23),
cout => N_52253,
dataf => N_52357,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_137\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_22_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_23\(34),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22.Z_CARRY_0\,
dataf => N_52365,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(334),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52251);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_22_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_80\(33),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22.Z_CARRY_1\,
dataf => N_52371,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_22\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_22_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_137\(32),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22.Z_CARRY_2\,
dataf => N_52372,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_79\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_22_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(22),
cout => N_52249,
dataf => N_52380,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_136\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_21_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_22\(35),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21.Z_CARRY_0\,
dataf => N_52388,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(333),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52247);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_21_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_79\(34),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21.Z_CARRY_1\,
dataf => N_52394,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_21\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_21_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_136\(33),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21.Z_CARRY_2\,
dataf => N_52395,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_78\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_21_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(21),
cout => N_52245,
dataf => N_52403,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_135\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_20_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_21\(36),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20.Z_CARRY_0\,
dataf => N_52411,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(332),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52243);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_20_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_78\(35),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20.Z_CARRY_1\,
dataf => N_52417,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_20\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_20_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_135\(34),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20.Z_CARRY_2\,
dataf => N_52418,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_77\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_20_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(20),
cout => N_52241,
dataf => N_52426,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_134\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_19_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_20\(37),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19.Z_CARRY_0\,
dataf => N_52434,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(331),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52239);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_19_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_77\(36),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19.Z_CARRY_1\,
dataf => N_52440,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_19\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_19_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_134\(35),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19.Z_CARRY_2\,
dataf => N_52441,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_76\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_19_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(19),
cout => N_52237,
dataf => N_52449,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_133\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_18_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_19\(38),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18.Z_CARRY_0\,
dataf => N_52457,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(330),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52235);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_18_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_76\(37),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18.Z_CARRY_1\,
dataf => N_52463,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_18\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_18_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_133\(36),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18.Z_CARRY_2\,
dataf => N_52464,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_75\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_18_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(18),
cout => N_52233,
dataf => N_52472,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_132\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_17_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_18\(39),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17.Z_CARRY_0\,
dataf => N_52480,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(329),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52231);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_17_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_75\(38),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17.Z_CARRY_1\,
dataf => N_52486,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_17\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_17_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_132\(37),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17.Z_CARRY_2\,
dataf => N_52487,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_74\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_17_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(17),
cout => N_52229,
dataf => N_52495,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_131\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_16_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_17\(40),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16.Z_CARRY_0\,
dataf => N_52503,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(328),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52227);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_16_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_74\(39),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16.Z_CARRY_1\,
dataf => N_52509,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_16\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_16_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_131\(38),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16.Z_CARRY_2\,
dataf => N_52510,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_73\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_16_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(16),
cout => N_52225,
dataf => N_52518,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_130\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_15_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_16\(41),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15.Z_CARRY_0\,
dataf => N_52526,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(327),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52223);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_15_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_73\(40),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15.Z_CARRY_1\,
dataf => N_52532,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_15\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_15_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_130\(39),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15.Z_CARRY_2\,
dataf => N_52533,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_72\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_15_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(15),
cout => N_52221,
dataf => N_52541,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_129\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_14_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_15\(42),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14.Z_CARRY_0\,
dataf => N_52549,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(326),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52219);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_14_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_72\(41),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14.Z_CARRY_1\,
dataf => N_52555,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_14\(43),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_14_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_129\(40),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14.Z_CARRY_2\,
dataf => N_52556,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_71\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_14_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(14),
cout => N_52217,
dataf => N_52564,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_128\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_13_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_14\(43),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13.Z_CARRY_0\,
dataf => N_52572,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(325),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52215);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_13_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_71\(42),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13.Z_CARRY_1\,
dataf => N_52578,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_13\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_13_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_128\(41),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13.Z_CARRY_2\,
dataf => N_52579,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_70\(43),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_13_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(13),
cout => N_52213,
dataf => N_52587,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_127\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_12_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_13\(44),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12.Z_CARRY_0\,
dataf => N_52595,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(324),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52211);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_12_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_70\(43),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12.Z_CARRY_1\,
dataf => N_52601,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_12\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_12_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_127\(42),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12.Z_CARRY_2\,
dataf => N_52602,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_69\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_12_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(12),
cout => N_52209,
dataf => N_52610,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_126\(43),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_11_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_12\(45),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11.Z_CARRY_0\,
dataf => N_52618,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(323),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52207);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_11_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_69\(44),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11.Z_CARRY_1\,
dataf => N_52624,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_11\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_11_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_126\(43),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11.Z_CARRY_2\,
dataf => N_52625,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_68\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_11_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(11),
cout => N_52205,
dataf => N_52633,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_125\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_10_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_11\(46),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10.Z_CARRY_0\,
dataf => N_52641,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(322),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52203);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_10_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_68\(45),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10.Z_CARRY_1\,
dataf => N_52647,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_10\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_10_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_125\(44),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10.Z_CARRY_2\,
dataf => N_52648,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_67\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_10_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(10),
cout => N_52201,
dataf => N_52656,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_124\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_39_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_40\(17),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39.Z_CARRY_0\,
dataf => N_52664,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(351),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_52199);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_39_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_97\(16),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39.Z_CARRY_1\,
dataf => N_52670,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_39\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_39_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_154\(15),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39.Z_CARRY_2\,
dataf => N_52671,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_96\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_39_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(39),
cout => N_52197,
dataf => N_52679,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_153\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_38_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_39\(18),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38.Z_CARRY_0\,
dataf => N_52687,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(350),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_52195);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_38_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_96\(17),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38.Z_CARRY_1\,
dataf => N_52693,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_38\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_38_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_153\(16),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38.Z_CARRY_2\,
dataf => N_52694,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_95\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_38_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(38),
cout => N_52193,
dataf => N_52702,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_152\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_37_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_38\(19),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37.Z_CARRY_0\,
dataf => N_52710,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(349),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_52191);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_37_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_95\(18),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37.Z_CARRY_1\,
dataf => N_52716,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_37\(20),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_37_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_152\(17),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37.Z_CARRY_2\,
dataf => N_52717,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_94\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_37_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(37),
cout => N_52189,
dataf => N_52725,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_151\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_36_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_37\(20),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36.Z_CARRY_0\,
dataf => N_52733,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(348),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_52187);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_36_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_94\(19),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36.Z_CARRY_1\,
dataf => N_52739,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_36\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_36_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_151\(18),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36.Z_CARRY_2\,
dataf => N_52740,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_93\(20),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_36_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(36),
cout => N_52185,
dataf => N_52748,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_150\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_35_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_36\(21),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35.Z_CARRY_0\,
dataf => N_52756,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(347),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_52183);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_35_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_93\(20),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35.Z_CARRY_1\,
dataf => N_52762,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_35\(22),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_35_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_150\(19),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35.Z_CARRY_2\,
dataf => N_52763,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_92\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_35_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(35),
cout => N_52181,
dataf => N_52771,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_149\(20),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_34_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_35\(22),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34.Z_CARRY_0\,
dataf => N_52779,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(346),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_52179);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_34_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_92\(21),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34.Z_CARRY_1\,
dataf => N_52785,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_34\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_34_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_149\(20),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34.Z_CARRY_2\,
dataf => N_52786,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_91\(22),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_34_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(34),
cout => N_52177,
dataf => N_52794,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_148\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_33_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_34\(23),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33.Z_CARRY_0\,
dataf => N_52802,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(345),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_52175);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_33_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_91\(22),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33.Z_CARRY_1\,
dataf => N_52808,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_33\(24),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_33_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_148\(21),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33.Z_CARRY_2\,
dataf => N_52809,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_90\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_33_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(33),
cout => N_52173,
dataf => N_52817,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_147\(22),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_32_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_33\(24),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32.Z_CARRY_0\,
dataf => N_52825,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(344),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_52171);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_32_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_90\(23),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32.Z_CARRY_1\,
dataf => N_52831,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_32\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_32_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_147\(22),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32.Z_CARRY_2\,
dataf => N_52832,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_89\(24),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_32_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(32),
cout => N_52169,
dataf => N_52840,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_146\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_31_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_32\(25),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31.Z_CARRY_0\,
dataf => N_52848,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(343),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52167);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_31_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_89\(24),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31.Z_CARRY_1\,
dataf => N_52854,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_31\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_31_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_146\(23),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31.Z_CARRY_2\,
dataf => N_52855,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_88\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_31_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(31),
cout => N_52165,
dataf => N_52863,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_145\(24),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_30_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_31\(26),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30.Z_CARRY_0\,
dataf => N_52871,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(342),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52163);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_30_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_88\(25),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30.Z_CARRY_1\,
dataf => N_52877,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_30\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_30_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_145\(24),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30.Z_CARRY_2\,
dataf => N_52878,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_87\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_30_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(30),
cout => N_52161,
dataf => N_52886,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_144\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_29_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_30\(27),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29.Z_CARRY_0\,
dataf => N_52894,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(341),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52159);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_29_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_87\(26),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29.Z_CARRY_1\,
dataf => N_52900,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_29\(28),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_29_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_144\(25),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29.Z_CARRY_2\,
dataf => N_52901,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_86\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_29_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(29),
cout => N_52157,
dataf => N_52909,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_143\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_28_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_29\(28),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28.Z_CARRY_0\,
dataf => N_52917,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(340),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52155);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_28_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_86\(27),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28.Z_CARRY_1\,
dataf => N_52923,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_28\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_28_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_143\(26),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28.Z_CARRY_2\,
dataf => N_52924,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_85\(28),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_28_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(28),
cout => N_52153,
dataf => N_52932,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_142\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_27_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_28\(29),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27.Z_CARRY_0\,
dataf => N_52940,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(339),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52151);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_27_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_85\(28),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27.Z_CARRY_1\,
dataf => N_52946,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_27\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_27_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_142\(27),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27.Z_CARRY_2\,
dataf => N_52947,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_84\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_27_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(27),
cout => N_52149,
dataf => N_52955,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_141\(28),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_26_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_27\(30),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26.Z_CARRY_0\,
dataf => N_52963,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(338),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52147);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_26_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_84\(29),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26.Z_CARRY_1\,
dataf => N_52969,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_26\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_26_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_141\(28),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26.Z_CARRY_2\,
dataf => N_52970,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_83\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_26_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(26),
cout => N_52145,
dataf => N_52978,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_140\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_25_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_26\(31),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25.Z_CARRY_0\,
dataf => N_52986,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(337),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52143);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_25_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_83\(30),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25.Z_CARRY_1\,
dataf => N_52992,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_25\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_25_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_140\(29),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25.Z_CARRY_2\,
dataf => N_52993,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_82\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_25_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(25),
cout => N_52141,
dataf => N_53001,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_139\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_5_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_6\(51),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5.Z_CARRY_0\,
dataf => N_53009,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(317),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52139);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_5_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_63\(50),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5.Z_CARRY_1\,
dataf => N_53015,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_5\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_5_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_120\(49),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5.Z_CARRY_2\,
dataf => N_53016,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_62\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_5_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(5),
cout => N_52137,
dataf => N_53024,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_119\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_4_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_5\(52),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4.Z_CARRY_0\,
dataf => N_53034,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(316),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52135);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_4_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000ff0")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_62\(51),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4.Z_CARRY_1\,
dataf => N_53044,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_12231\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5771\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_4_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000ff0")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_119\(50),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4.Z_CARRY_2\,
dataf => N_53045,
datad => N_30731,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6583\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_4_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000ff0")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(4),
cout => N_52133,
dataf => N_53049,
datad => N_53048,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_60\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6961\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_52_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_53\(4),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52.Z_CARRY_0\,
dataf => N_53054,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(364),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_52131);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_52_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_110\(3),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52.Z_CARRY_1\,
dataf => N_53060,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_52\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_52_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_167\(2),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52.Z_CARRY_2\,
dataf => N_53061,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_109\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_52_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(52),
cout => N_52129,
dataf => N_53069,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_166\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_51_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_52\(5),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51.Z_CARRY_0\,
dataf => N_53077,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(363),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_52127);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_51_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_109\(4),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51.Z_CARRY_1\,
dataf => N_53083,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_51\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_51_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_166\(3),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51.Z_CARRY_2\,
dataf => N_53084,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_108\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_51_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(51),
cout => N_52125,
dataf => N_53092,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_165\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_50_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_51\(6),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50.Z_CARRY_0\,
dataf => N_53100,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(362),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_52123);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_50_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_108\(5),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50.Z_CARRY_1\,
dataf => N_53106,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_50\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_50_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_165\(4),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50.Z_CARRY_2\,
dataf => N_53107,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_107\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_50_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(50),
cout => N_52121,
dataf => N_53115,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_164\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_49_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_50\(7),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49.Z_CARRY_0\,
dataf => N_53123,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(361),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_52119);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_49_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_107\(6),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49.Z_CARRY_1\,
dataf => N_53129,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_49\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_49_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_164\(5),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49.Z_CARRY_2\,
dataf => N_53130,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_106\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_49_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(49),
cout => N_52117,
dataf => N_53138,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_163\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_48_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_49\(8),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48.Z_CARRY_0\,
dataf => N_53146,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(360),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_52115);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_48_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_106\(7),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48.Z_CARRY_1\,
dataf => N_53152,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_48\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_48_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_163\(6),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48.Z_CARRY_2\,
dataf => N_53153,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_105\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_48_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(48),
cout => N_52113,
dataf => N_53161,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_162\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_47_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_48\(9),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47.Z_CARRY_0\,
dataf => N_53169,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(359),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_52111);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_47_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_105\(8),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47.Z_CARRY_1\,
dataf => N_53175,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_47\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_47_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_162\(7),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47.Z_CARRY_2\,
dataf => N_53176,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_104\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_47_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(47),
cout => N_52109,
dataf => N_53184,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_161\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_46_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_47\(10),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46.Z_CARRY_0\,
dataf => N_53192,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(358),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_52107);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_46_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_104\(9),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46.Z_CARRY_1\,
dataf => N_53198,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_46\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_46_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_161\(8),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46.Z_CARRY_2\,
dataf => N_53199,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_103\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_46_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(46),
cout => N_52105,
dataf => N_53207,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_160\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_45_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_46\(11),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45.Z_CARRY_0\,
dataf => N_53215,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(357),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_52103);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_45_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_103\(10),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45.Z_CARRY_1\,
dataf => N_53221,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_45\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_45_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_160\(9),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45.Z_CARRY_2\,
dataf => N_53222,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_102\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_45_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(45),
cout => N_52101,
dataf => N_53230,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_159\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_44_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_45\(12),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44.Z_CARRY_0\,
dataf => N_53238,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(356),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_52099);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_44_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_102\(11),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44.Z_CARRY_1\,
dataf => N_53244,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_44\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_44_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_159\(10),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44.Z_CARRY_2\,
dataf => N_53245,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_101\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_44_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(44),
cout => N_52097,
dataf => N_53253,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_158\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_43_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_44\(13),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43.Z_CARRY_0\,
dataf => N_53261,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(355),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_52095);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_43_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_101\(12),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43.Z_CARRY_1\,
dataf => N_53267,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_43\(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_43_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_158\(11),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43.Z_CARRY_2\,
dataf => N_53268,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_100\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_43_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(43),
cout => N_52093,
dataf => N_53276,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_157\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_42_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_43\(14),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42.Z_CARRY_0\,
dataf => N_53284,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(354),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_52091);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_42_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_100\(13),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42.Z_CARRY_1\,
dataf => N_53290,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_42\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_42_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_157\(12),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42.Z_CARRY_2\,
dataf => N_53291,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_99\(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_42_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(42),
cout => N_52089,
dataf => N_53299,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_156\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_41_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_42\(15),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41.Z_CARRY_0\,
dataf => N_53307,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(353),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_52087);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_41_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_99\(14),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41.Z_CARRY_1\,
dataf => N_53313,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_41\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_41_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_156\(13),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41.Z_CARRY_2\,
dataf => N_53314,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_98\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_41_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(41),
cout => N_52085,
dataf => N_53322,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_155\(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_40_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_41\(16),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40.Z_CARRY_0\,
dataf => N_53330,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(352),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_52083);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_40_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_98\(15),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40.Z_CARRY_1\,
dataf => N_53336,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_40\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_40_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_155\(14),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40.Z_CARRY_2\,
dataf => N_53337,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_97\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_40_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(40),
cout => N_52081,
dataf => N_53345,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_154\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff0000f0cc")
port map (
sumout => \GRLFPC2_0.FPO.EXP\(0),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10870\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10857\,
cin => N_52079);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff0000f3c0")
port map (
sumout => \GRLFPC2_0.FPO.EXP\(1),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10858\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10871\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff0000f3c0")
port map (
sumout => \GRLFPC2_0.FPO.EXP\(2),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10859\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10872\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff0000f3c0")
port map (
sumout => \GRLFPC2_0.FPO.EXP\(3),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10860\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10873\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_4: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff0000f3c0")
port map (
sumout => \GRLFPC2_0.FPO.EXP\(4),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10861\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10874\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_5: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff0000fc30")
port map (
sumout => \GRLFPC2_0.FPO.EXP\(5),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10875\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10862\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_4\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_6: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff0000fc30")
port map (
sumout => \GRLFPC2_0.FPO.EXP\(6),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10876\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10862\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_5\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_7: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff0000fc30")
port map (
sumout => \GRLFPC2_0.FPO.EXP\(7),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10877\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10864\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_6\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_8: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff0000fc30")
port map (
sumout => \GRLFPC2_0.FPO.EXP\(8),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10878\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10864\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_7\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_9: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff0000f3c0")
port map (
sumout => \GRLFPC2_0.FPO.EXP\(9),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_9\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10864\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10879\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_8\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_10: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cc330000f000")
port map (
sumout => \GRLFPC2_0.FPO.EXP\(10),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_10\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5301\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10880\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_9\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_11: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cc330000f000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(11),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_11\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5343\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10881\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_10\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_12: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cc330000f000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(12),
cout => N_8,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5339\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10882\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_11\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_3_0_RNIRC7P: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ccff0000f000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_57\(0),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(368),
datad => N_53417,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
cin => N_52075);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_0_RNI7BMN1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00003000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SBLSBS_1\(1),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_56\(1),
datad => N_53423,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_1_0_RNICAOM3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SCLSBS_2\(0),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_2\,
dataf => N_53424,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_113\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_1_0_RNICAOM3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_954\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_3\,
dataf => VCC,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_1_0_RNI0DGF7: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN25_NOTPROP\,
cout => N_52073,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SCLSBS_1\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_55_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_56\(1),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55.Z_CARRY_0\,
dataf => N_53435,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(367),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_52071);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_55_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_113\(0),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55.Z_CARRY_1\,
dataf => N_53441,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_55\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_55_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SCLSBS_1\(1),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55.Z_CARRY_2\,
dataf => N_53442,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_112\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_55_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000c00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(55),
cout => N_52069,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI\(0),
datad => N_53450,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_54_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_55\(2),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54.Z_CARRY_0\,
dataf => N_53458,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(366),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_52067);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_54_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_112\(1),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54.Z_CARRY_1\,
dataf => N_53464,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_54\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_54_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI\(0),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54.Z_CARRY_2\,
dataf => N_53465,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_111\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_54_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(54),
cout => N_52065,
dataf => N_53473,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_168\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_53_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_54\(3),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53.Z_CARRY_0\,
dataf => N_53481,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(365),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
cin => N_52063);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_53_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_111\(2),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53.Z_CARRY_1\,
dataf => N_53487,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_53\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_53_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_168\(1),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53.Z_CARRY_2\,
dataf => N_53488,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_110\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_53_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(53),
cout => N_52061,
dataf => N_53496,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_167\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_7_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_8\(49),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7.Z_CARRY_0\,
dataf => N_53504,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(319),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52059);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_7_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_65\(48),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7.Z_CARRY_1\,
dataf => N_53510,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_7\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_7_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_122\(47),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7.Z_CARRY_2\,
dataf => N_53511,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_64\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_7_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(7),
cout => N_52057,
dataf => N_53519,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_121\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_6_Z_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000033ff00000f00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_7\(50),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6.Z_CARRY_0\,
dataf => N_53527,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(318),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
cin => N_52055);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_6_Z_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_64\(49),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6.Z_CARRY_1\,
dataf => N_53533,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_6\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6.Z_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_6_Z_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cfff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_121\(48),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6.Z_CARRY_2\,
dataf => N_53534,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_63\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6.Z_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_6_Z_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3ff0000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(6),
cout => N_52053,
dataf => N_53542,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_120\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6.Z_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_6_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(63),
cout => N_9,
cin => N_52053);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_6_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52055,
datad => N_53526,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_7_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(64),
cin => N_52057);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_7_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52059,
datad => N_53503,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_53_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(110),
cin => N_52061);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_53_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52063,
datad => N_53480,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_54_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(111),
cin => N_52065);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_54_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52067,
datad => N_53457,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_55_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(112),
cin => N_52069);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_55_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52071,
datad => N_53434,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN2_MIXOIN_3_RNO_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_4\,
cin => N_52073);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_RNIUKAC_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52075,
datad => N_53416,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000f0cc")
port map (
cout => N_52079,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_40_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(97),
cin => N_52081);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_40_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52083,
datad => N_53329,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_41_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(98),
cin => N_52085);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_41_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52087,
datad => N_53306,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_42_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(99),
cin => N_52089);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_42_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52091,
datad => N_53283,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_43_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(100),
cin => N_52093);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_43_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52095,
datad => N_53260,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_44_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(101),
cin => N_52097);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_44_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52099,
datad => N_53237,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_45_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(102),
cin => N_52101);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_45_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52103,
datad => N_53214,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_46_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(103),
cin => N_52105);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_46_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52107,
datad => N_53191,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_47_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(104),
cin => N_52109);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_47_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52111,
datad => N_53168,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_48_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(105),
cin => N_52113);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_48_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52115,
datad => N_53145,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_49_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(106),
cin => N_52117);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_49_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52119,
datad => N_53122,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_50_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(107),
cin => N_52121);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_50_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52123,
datad => N_53099,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_51_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(108),
cin => N_52125);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_51_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52127,
datad => N_53076,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_52_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(109),
cin => N_52129);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_52_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52131,
datad => N_53053,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_4_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(61),
cin => N_52133);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_4_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52135,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10626\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_5_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(62),
cin => N_52137);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_5_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52139,
datad => N_53008,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_25_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(82),
cin => N_52141);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_25_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52143,
datad => N_52985,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_26_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(83),
cin => N_52145);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_26_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52147,
datad => N_52962,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_27_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(84),
cin => N_52149);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_27_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52151,
datad => N_52939,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_28_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(85),
cin => N_52153);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_28_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52155,
datad => N_52916,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_29_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(86),
cin => N_52157);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_29_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52159,
datad => N_52893,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_30_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(87),
cin => N_52161);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_30_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52163,
datad => N_52870,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_31_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(88),
cin => N_52165);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_31_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52167,
datad => N_52847,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_32_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(89),
cin => N_52169);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_32_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52171,
datad => N_52824,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_33_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(90),
cin => N_52173);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_33_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52175,
datad => N_52801,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_34_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(91),
cin => N_52177);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_34_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52179,
datad => N_52778,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_35_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(92),
cin => N_52181);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_35_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52183,
datad => N_52755,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_36_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(93),
cin => N_52185);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_36_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52187,
datad => N_52732,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_37_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(94),
cin => N_52189);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_37_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52191,
datad => N_52709,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_38_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(95),
cin => N_52193);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_38_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52195,
datad => N_52686,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_39_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(96),
cin => N_52197);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_39_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52199,
datad => N_52663,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_10_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(67),
cin => N_52201);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_10_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52203,
datad => N_52640,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_11_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(68),
cin => N_52205);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_11_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52207,
datad => N_52617,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_12_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(69),
cin => N_52209);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_12_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52211,
datad => N_52594,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_13_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(70),
cin => N_52213);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_13_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52215,
datad => N_52571,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_14_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(71),
cin => N_52217);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_14_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52219,
datad => N_52548,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_15_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(72),
cin => N_52221);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_15_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52223,
datad => N_52525,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_16_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(73),
cin => N_52225);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_16_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52227,
datad => N_52502,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_17_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(74),
cin => N_52229);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_17_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52231,
datad => N_52479,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_18_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(75),
cin => N_52233);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_18_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52235,
datad => N_52456,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_19_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(76),
cin => N_52237);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_19_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52239,
datad => N_52433,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_20_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(77),
cin => N_52241);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_20_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52243,
datad => N_52410,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_21_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(78),
cin => N_52245);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_21_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52247,
datad => N_52387,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_22_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(79),
cin => N_52249);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_22_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52251,
datad => N_52364,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_23_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(80),
cin => N_52253);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_23_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52255,
datad => N_52341,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_24_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(81),
cin => N_52257);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_24_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52259,
datad => N_52318,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_8_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(65),
cin => N_52261);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_8_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52263,
datad => N_52295,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_9_Z_CARRY_3_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(66),
cin => N_52265);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_9_Z_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000cf00")
port map (
cout => N_52267,
datad => N_52272,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
cin => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_0_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"cfc0ffff8a80a0a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_0_0_13__G0_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(13),
datae => \GRLFPC2_0.FPI.LDOP_0_0\,
datad => N_633,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3639\,
datab => N_697,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4534\,
datag => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_1_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"d0d0dd0dd0d00d0d")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_1\(0),
dataf => \GRLFPC2_0.R.I.EXC\(0),
datae => \GRLFPC2_0.N_1517\,
datad => \GRLFPC2_0.R.FSR.TEM\(0),
datac => \GRLFPC2_0.N_1015\,
datab => N_366,
dataa => \GRLFPC2_0.V.FSR.CEXC_2_SQMUXA\,
datag => N_406);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_1_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"d0d0dd0dd0d00d0d")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_1\(2),
dataf => \GRLFPC2_0.R.I.EXC\(2),
datae => \GRLFPC2_0.N_1517\,
datad => \GRLFPC2_0.R.FSR.TEM\(2),
datac => \GRLFPC2_0.N_1015\,
datab => N_368,
dataa => \GRLFPC2_0.V.FSR.CEXC_2_SQMUXA\,
datag => N_408);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_10: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"faf5f9f9af5f9f9f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_10\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10871\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10857\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10858\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(1),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10870\);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_1_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"d0d0dd0dd0d00d0d")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_1\(1),
dataf => \GRLFPC2_0.R.I.EXC\(1),
datae => \GRLFPC2_0.N_1517\,
datad => \GRLFPC2_0.R.FSR.TEM\(1),
datac => \GRLFPC2_0.N_1015\,
datab => N_367,
dataa => \GRLFPC2_0.V.FSR.CEXC_2_SQMUXA\,
datag => N_407);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_1_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"d0d0dd0dd0d00d0d")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_1\(3),
dataf => \GRLFPC2_0.R.I.EXC\(3),
datae => \GRLFPC2_0.N_1517\,
datad => \GRLFPC2_0.R.FSR.TEM\(3),
datac => \GRLFPC2_0.N_1015\,
datab => N_369,
dataa => \GRLFPC2_0.V.FSR.CEXC_2_SQMUXA\,
datag => N_409);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_1_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"d0d0dd0dd0d00d0d")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_1\(4),
dataf => \GRLFPC2_0.R.I.EXC\(4),
datae => \GRLFPC2_0.N_1517\,
datad => \GRLFPC2_0.R.FSR.TEM\(4),
datac => \GRLFPC2_0.N_1015\,
datab => N_370,
dataa => \GRLFPC2_0.V.FSR.CEXC_2_SQMUXA\,
datag => N_410);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_234_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"b3a0b3a0a0a0a0a0")
port map (
combout => N_37230,
dataf => \GRLFPC2_0.FPI.LDOP_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datad => \GRLFPC2_0.FPI.OP2\(62),
datac => \GRLFPC2_0.FPO.EXP\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
dataa => N_37019_2,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(247));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_235_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"b3a0b3a0a0a0a0a0")
port map (
combout => N_37203,
dataf => \GRLFPC2_0.FPI.LDOP_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datad => \GRLFPC2_0.FPI.OP2\(61),
datac => \GRLFPC2_0.FPO.EXP\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
dataa => N_37019_2,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_236_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"b3a0b3a0a0a0a0a0")
port map (
combout => N_37176,
dataf => \GRLFPC2_0.FPI.LDOP_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datad => \GRLFPC2_0.FPI.OP2\(60),
datac => \GRLFPC2_0.FPO.EXP\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
dataa => N_37019_2,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(249));
\GRLFPC2_0_COMB_RF2REN_1_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"4477747444747474")
port map (
combout => RFI2_REN2Z,
dataf => \GRLFPC2_0.COMB.RS2_1\(0),
datae => N_13,
datad => \GRLFPC2_0.N_3477_1_I\,
datac => \GRLFPC2_0.R.A.RF2REN\(2),
datab => N_398,
dataa => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT\,
datag => \GRLFPC2_0.COMB.RS2D_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"fe54f5f5fe54a0a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f00ff00f88778877")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(226),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f00ff00f88778877")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(31),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(200),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_30_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f00ff00f88778877")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(30),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(201),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f00ff00f88778877")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(228),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f00ff00f88778877")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(8),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(223),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f00ff00f88778877")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(33),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(198),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_35_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f00ff00f88778877")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(35),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(196),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"9a95a5a59a955555")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(49),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(182),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f00ff00f88778877")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(225),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f00ff00f88778877")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(32),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(199),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_37_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f00ff00f88778877")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(37),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(194),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"9a95a5a59a955555")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(24),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(207),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f00ff00f88778877")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(224),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_9_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(9),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(222),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_16_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(16),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(215),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(36),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(195),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(28),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(203),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(178),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_23_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(23),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(208),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_15_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(15),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(216),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(184),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(177),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(17),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(214),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(48),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(183),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(18),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(213),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(39),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(192),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_22_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(22),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(209),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(176),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(50),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(181),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_41_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(41),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(190),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"5565669555655595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(29),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(202),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5346\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(12),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(219),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(34),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(197),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(56),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(175),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_40_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(40),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(191),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_44_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(44),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(187),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(52),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(179),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(13),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(218),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(27),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(204),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_46_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(46),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(185),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(19),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(212),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_20_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(20),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(211),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(38),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(193),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"ff008080f0008080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_1\,
dataf => N_32844_3,
datae => N_29071_1,
datad => N_32723_1,
datac => N_32861_1,
datab => N_33140_1,
dataa => N_32730_1,
datag => N_33340_I);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_43_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(43),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(188),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(42),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(189),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(26),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(205),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(11),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(220),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(25),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(206),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(51),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(180),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_14_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(14),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(217),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_21_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(21),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(210),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"a5aa9595a5559595")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(10),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(221),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_2_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"3000120000000000")
port map (
combout => N_34257,
dataf => N_29195_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81),
datag => N_33436_1);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f6f9f9f96f9f9f9f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10881\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10861\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5343\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10874\);
GRLFPC2_0_COMB_ANNULRES_1_IV_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"fff0f8f8fff00808")
port map (
combout => \GRLFPC2_0.N_82\,
dataf => \GRLFPC2_0.N_1683\,
datae => \GRLFPC2_0.R.M.FPOP\,
datad => N_295,
datac => \GRLFPC2_0.R.E.FPOP\,
datab => \GRLFPC2_0.N_1685\,
dataa => \GRLFPC2_0.R.A.FPOP\,
datag => N_294);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_0_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"efefdecfffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_0\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83),
datag => N_32844_3);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"000f404000004040")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_0\,
dataf => N_28211_1,
datae => N_34029,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_604\,
datac => N_28892_I,
datab => N_33503_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_7_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"afffffffaeeeefef")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_7\(11),
dataf => N_33055,
datae => N_32730_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78),
datac => N_32959_I,
datab => N_33179,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_1_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"0000000004000400")
port map (
combout => N_34182,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_531\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"e0eee0ee00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_1\,
datae => N_27258,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\,
datac => N_27315,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
datag => N_27316);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIK8286_20_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f0f00000f0f0fd02")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datae => \GRLFPC2_0.FPI.LDOP_0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(20),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11));
GRLFPC2_0_COMB_RDD_1_M11: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"0500000000000020")
port map (
combout => \GRLFPC2_0.COMB.RDD_1.N_12\,
dataf => N_72,
datae => N_73,
datad => N_83,
datac => \GRLFPC2_0.N_624_3\,
datab => \GRLFPC2_0.COMB.RDD_1.N_27\,
dataa => N_76,
datag => N_74);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_1_A3_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"1555505015555555")
port map (
combout => N_28510,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1636\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(249),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_I_O2_3_0\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1637\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(247));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN20_LOCOV: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"fffeeaeafffaaaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5330\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.REEXCOVUV.UN13_LOCOV_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\,
datad => \GRLFPC2_0.FPO.EXP\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5335\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.REEXCOVUV.UN13_LOCOV_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(11),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.REEXCOVUV.UN25_LOCOV_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"000a808000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_12\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82),
datac => N_33607_1,
datab => N_33984_2,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85),
datag => N_33111);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_9_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"0050010100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_5\,
dataf => N_28271_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_782\,
datab => N_32979_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_604\,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_603\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_0_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"ffffffeff33fffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_0\(60),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datad => N_34239_I,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_24_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"0000000002000200")
port map (
combout => N_32902,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_603\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_0_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"0208020800000000")
port map (
combout => N_34181,
dataf => N_33659_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M12_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f0fff2f2f0f0f2f2")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7350\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M12_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"0f0f0e0e0f000e0e")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7350\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M13_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f0fff2f2f0f0f2f2")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7352\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_YY_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"0000323200033232")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7778\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7352\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM6\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_24_RNI32HA1_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"3bffb1f5ce0ae4a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO5_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_8\,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_30_RNI02HA1_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"3bffb1f5ce0ae4a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_8\,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_12: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(12),
cout => N_10,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(232),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(245),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_11\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_11: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(11),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_11\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_10\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_10: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(10),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_10\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(247),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_9\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_9: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(9),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_9\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_8\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_8: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(8),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(249),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_7\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_7: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(7),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(237),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(250),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_6\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_6: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(6),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(238),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(251),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_5\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_5: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(5),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(239),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(252),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_4\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_4: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(4),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(240),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(253),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(3),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(241),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(254),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(2),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(255),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(1),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(256),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000ff00")
port map (
sumout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(0),
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(257),
cin => N_66927);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CARRY_0_BUF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ff00")
port map (
cout => N_66927,
datad => VCC,
cin => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffbfffff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7248\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_0_0_13__G0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4534\,
datad => \GRLFPC2_0.FPI.LDOP_0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12));
GRLFPC2_0_COMB_V_MK_BUSY_2_I_O3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffdfffffffffff")
port map (
combout => \GRLFPC2_0.N_3545\,
dataf => \GRLFPC2_0.FPO.BUSY_O\,
datae => \GRLFPC2_0.R.MK.RST_O_0\,
datad => \GRLFPC2_0.R.MK.HOLDN2_O_0\,
datac => \GRLFPC2_0.R.MK.HOLDN1_O_0\,
datab => \GRLFPC2_0.R.MK.RST2_O_0\,
dataa => RST_RETO);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffca0000ff35")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_I_I_0\(0),
datae => N_66617,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP\,
datab => N_36985,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_0_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff0f33ffff")
port map (
combout => N_66617,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP\,
datac => N_36986,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0cc00000f33")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4424\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_I_I_0\(0),
datae => N_66615,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP\,
datac => N_36985,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_0_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff0f0fffffffff")
port map (
combout => N_66615,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP\,
datad => N_36986,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_7_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000c000c333f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_3_RETI\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10066\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10067\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10126\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10127\,
datab => N_61587_I_0);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_4_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3fff3fff3ccc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM6_RETI\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10067\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10066\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10127\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10126\,
datab => N_61587_I_0);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_RNI1ET3Q22_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff0ff707")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_6__G2\,
dataf => N_66607,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10128\,
datac => N_61587_I_0,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIM9ICH22_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0004003400070037")
port map (
combout => N_66607,
dataf => \GRLFPC2_0.FPO.FRAC\(51),
datae => \GRLFPC2_0.FPO.FRAC\(50),
datad => N_61587_I_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_RNIT582FG2_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff0ff707")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_11__G2\,
dataf => N_66597,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10123\,
datac => N_61587_I_0,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNI82VQ5G2_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0004003400070037")
port map (
combout => N_66597,
dataf => \GRLFPC2_0.FPO.FRAC\(46),
datae => \GRLFPC2_0.FPO.FRAC\(45),
datad => N_61587_I_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIJQBD1U1_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fffe0000f7f6")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_12__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(12),
datae => N_66595,
datad => \GRLFPC2_0.FPO.FRAC\(45),
datac => N_61587_I_0,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_RNI8IEMPR_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0004ff040034ff34")
port map (
combout => N_66595,
dataf => \GRLFPC2_0.FPO.FRAC\(44),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10122\,
datad => N_61587_I_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_RNISETO9G1_14_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff0ff707")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_14__G2\,
dataf => N_66593,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(14),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10120\,
datac => N_61587_I_0,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNILPF90G1_15_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0004003400070037")
port map (
combout => N_66593,
dataf => \GRLFPC2_0.FPO.FRAC\(43),
datae => \GRLFPC2_0.FPO.FRAC\(42),
datad => N_61587_I_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIPNQN9C_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fffe0000f7f6")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_17__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(17),
datae => N_66587,
datad => \GRLFPC2_0.FPO.FRAC\(40),
datac => N_61587_I_0,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_RNIA62NTL1_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0004ff040034ff34")
port map (
combout => N_66587,
dataf => \GRLFPC2_0.FPO.FRAC\(39),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10117\,
datad => N_61587_I_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNINAR1SC3_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fffe0000f7f6")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_16__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(16),
datae => N_66585,
datad => \GRLFPC2_0.FPO.FRAC\(41),
datac => N_61587_I_0,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_RNI8D3P3M2_16_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0004ff040034ff34")
port map (
combout => N_66585,
dataf => \GRLFPC2_0.FPO.FRAC\(40),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10118\,
datad => N_61587_I_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNI0DGN0E1_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fffb0000f7f3")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_15__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(15),
datae => N_66583,
datad => \GRLFPC2_0.FPO.FRAC\(41),
datac => N_61587_I_0,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_RNIMVB58N_15_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0004ff040007ff07")
port map (
combout => N_66583,
dataf => \GRLFPC2_0.FPO.FRAC\(42),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10119\,
datad => N_61587_I_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_RNIQBNIKU1_9_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff0ff707")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_9__G2\,
dataf => N_66581,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10125\,
datac => N_61587_I_0,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNI0RN2BU1_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0004003400070037")
port map (
combout => N_66581,
dataf => \GRLFPC2_0.FPO.FRAC\(48),
datae => \GRLFPC2_0.FPO.FRAC\(47),
datad => N_61587_I_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fff3000033f3")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
dataf => N_27316,
datae => N_66571,
datad => N_27258,
datac => N_27315,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_SUB: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000003ffffffff")
port map (
combout => N_66571,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_1\,
datae => \GRLFPC2_0.FPI.LDOP_0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_RNO_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff00fe00fb00fa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_1__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_176__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_175__G2\,
datad => N_66569,
datac => N_61587_I_0,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_RNO_0_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000400c4ff04ffc4")
port map (
combout => N_66569,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10133\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(1),
datad => N_61587_I_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_2_IV_RNO_0_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"5555050105010501")
port map (
combout => N_65541,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_49_I\,
datac => \GRLFPC2_0.FPI.LDOP_0_0\,
datab => N_66565,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_2_IV_RNO_1_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000fffffff0")
port map (
combout => N_66565,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4238\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_17_RNO_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000023f300002fff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_386\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN11_WQSTSETS\,
datae => N_66563,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_17_RNO_0_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fff0fff0fff0")
port map (
combout => N_66563,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1677\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1770\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_547\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233));
GRLFPC2_0_R_MK_BUSY_RET_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffff3fcfcfcf0")
port map (
combout => \GRLFPC2_0.R.MK.BUSY_RET_0_0_G0_MUX2\,
dataf => D_N_7,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\,
datad => N_65488,
datac => N_65602,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M5S4: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffd8")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7350_RETI\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_11__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_12__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_14__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10061\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10121\,
dataa => N_61587_I_0);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M5_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000c3f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5_RETI\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_11__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_12__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10061\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10121\,
datab => N_61587_I_0);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_1_RNIBRMR: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0dcddfdff2322020")
port map (
combout => N_30731,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10626\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(316));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_12_RNI97FJ5_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"5555555544440040")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_49_I\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1544\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1852\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1503\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1633\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1618\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN5_ZERO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33ff5f5fffccfafa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_6_RNI66SI: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0000000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(109),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_RETO\,
datad => \GRLFPC2_0.FPI.LDOP_I_RETO\,
datac => RFO2_DATA1_RETO(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_1_RNI02SI: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0000000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(108),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_RETO\,
datad => \GRLFPC2_0.FPI.LDOP_I_RETO\,
datac => RFO2_DATA1_RETO(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_0__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10074\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10134\,
datad => N_61587_I_0);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_66446,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_0__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_66445,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_2__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_66444,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_4__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_0_C: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00c00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_TZ\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_513\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1809\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_479\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_141_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(141),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_14\(141),
datae => \GRLFPC2_0.FPO.FRAC\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_31_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1770\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(249),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(247));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPYBUS_2_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPYBUS_2_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_30_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1677\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_O2_10_4_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_O2_10_4\(83),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(253),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(251),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(257),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(252));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_80_RNI0SCO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1637\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(250),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(255),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(254),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(253),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_I_O2_4_4\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_115_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000c000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(115),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(118));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_71_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(71),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datae => N_27258,
datad => N_27290,
datac => N_27289,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_71_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccccccff00f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(71),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datae => N_27258,
datad => N_27286,
datac => N_27285,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_M2_E_RNI5AEF943: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0f0f030c0c0c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M\(3),
dataf => D_N_7,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\,
datad => N_65488,
datac => N_65578,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_M2_E_RNIPAOD943: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0f0f030c0c0c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M\(1),
dataf => D_N_7,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\,
datad => N_65488,
datac => N_65584,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_0_D: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f4f1f1f1f5")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D\,
dataf => D_N_7,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\,
datad => N_65488,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_90_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cccccc4e8d8d8d0f")
port map (
combout => N_65609,
dataf => D_N_7,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\,
datad => N_65488,
datac => N_65588,
datab => N_65572,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_M2_E_RNIGA3K253: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000080404040c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1\,
dataf => D_N_7,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\,
datad => N_65488,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_51_I\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_PCTRL_NEW_1_S_RNIBDU7943: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333333b3737373f3")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1\,
dataf => D_N_7,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\,
datad => N_65488,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_O2_11_3_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ffffffffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_O2_11_3\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(237));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_72_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(72),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(43),
datac => \GRLFPC2_0.FPO.FRAC\(41),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaff00f0f0cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(60),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_176__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaff00f0f0cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(59),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_175__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_M2_E_RNI0VH3C43: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffff3fcfcfcf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0\,
dataf => D_N_7,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\,
datad => N_65488,
datac => N_65570,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_PCTRL_NEW_1_S_RNI43MGH43: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c3c003c003c003c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_N_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_N_4\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_0_0_TZ_RNIFG4K843: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000004010101050")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0\,
dataf => D_N_7,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\,
datad => N_65488,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_TZ\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIELMI_231_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.EXTEND.TEMP_0\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5346\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(15),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(231));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_84_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(84),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_85_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(85),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_86_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(86),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(86),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(86),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_105_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(105),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(105),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(105),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_104_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(104),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(104),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(104),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_102_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(102),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(102),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(102),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_80_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_79_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_100_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(100),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(100),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(100),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_64_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(64),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(64),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(64),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_99_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(99),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(99),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(99),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_98_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(98),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(98),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(98),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_97_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(97),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(97),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(97),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_89_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(89),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(89),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(89));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_87_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(87),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(87),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(87),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_88_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(88),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(88),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(88));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_96_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(96),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(96),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(96),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_90_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(90),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(90),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(90));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_95_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(95),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(95),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(95),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_77_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(77),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(77),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(77),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_92_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(92),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(92),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(92),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_94_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(94),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(94),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(94),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_76_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(76),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(76),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(76),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_74_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(74),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(74),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(74),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_141_RNIEGLM: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
dataf => \GRLFPC2_0.FPI.LDOP_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(80));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_138_RNIQ8LM: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
dataf => \GRLFPC2_0.FPI.LDOP_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_72_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(72),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(72),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(72));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_130_RNI1EO51: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(115),
dataf => \GRLFPC2_0.FPI.LDOP_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1_RETO\(115),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0_RETO\(115));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_127_RNIM0LM: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
dataf => \GRLFPC2_0.FPI.LDOP_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(64),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(64));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_124_RNIG0LM: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
dataf => \GRLFPC2_0.FPI.LDOP_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(77),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(77));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_121_RNIA0LM: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
dataf => \GRLFPC2_0.FPI.LDOP_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(76),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(76));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_118_RNIMOKM: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
dataf => \GRLFPC2_0.FPI.LDOP_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(74),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(74));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_RNI7DIK_72_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(72),
datae => \GRLFPC2_0.FPI.LDOP_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(72));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_71_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccccccff00f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(71),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1_RETO\(71),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0_RETO\(71),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(71));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_RNI79IK_71_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(71),
datae => \GRLFPC2_0.FPI.LDOP_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(71));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_400_RNIBQ6O: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datae => N_65488_RETO_0,
datad => D_N_7_RETO_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_102_RNIQ1N51: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000cc000000f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO\,
datae => \GRLFPC2_0.FPI.LDOP_1_RETO\,
datad => \GRLFPC2_0.FPI.RST_1_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(113),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_372__G1_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_SUB_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc0fffffcc0fff")
port map (
combout => N_65516,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(43));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_97_RNIJVT21: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffccfffffff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO\,
datae => \GRLFPC2_0.FPI.LDOP_1_RETO\,
datad => \GRLFPC2_0.FPI.RST_1_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_319__G1_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPYBUS_2_9_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2_RETI\(9),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(29),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(30),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_80_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fffffffffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_I_O2_4_4_RETI\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(251),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(252),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(256),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(257));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNI8OPN_227_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10746\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5346\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(227));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIAOPN_229_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10744\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5346\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(229));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_92_RNI9VT21: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000cc000000f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO\,
datae => \GRLFPC2_0.FPI.LDOP_1_RETO\,
datad => \GRLFPC2_0.FPI.RST_1_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_318__G1_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_109_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccff00f0f0ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(109),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_RETO\,
datae => N_58999_RETO,
datad => N_59000_RETO,
datac => \GRLFPC2_0.FPO.FRAC_RETO\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_108_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccff00f0f0ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(108),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_RETO\,
datae => N_58999_RETO,
datad => N_59001_RETO,
datac => \GRLFPC2_0.FPO.FRAC_RETO\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(50));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_76_RNI7D391: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000aaaaf0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114),
dataf => \GRLFPC2_0.FPI.LDOP_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1_RETO\(114),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0_RETO\(114),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_3_I_RETO\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_90_RNI0RBU: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fff00ff00ff00ff")
port map (
combout => N_65771_RETO,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO\,
datad => N_65609_RETO,
datac => CPI_D_INST_RETO(7));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_74_RNIB3U21: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c3cff3caa3caa3c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO5_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_65_RNIG1E21_5: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333030033330000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_TZ_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datab => CPI_D_INST_RETO(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_28_RNIJ1E21_7: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c333003300330033")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(84));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_55_RNIR4BR_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff0fff0ccf0ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000300f300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_9\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_30_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(30),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_30__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(29),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_COMPUTECONST_UN25_RESVEC: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC_RETI\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(29),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(30),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_43_RNIEOHD1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffefffcfffcfffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO\,
dataa => CPI_D_INST_RETO(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_YY_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000afae00000504")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7786\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M11\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7352\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M11_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffffff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M11\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_COUNTSUCCESSIVEZERO36_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_0_RETI\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_6__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_16__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(12),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNI9GTI_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ff00f0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5346_RETI\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(374),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_XX_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000bbbbbbb8")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7777\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7350\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M14S2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM12\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7352\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_7__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10067\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10127\,
datad => N_61587_I_0);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_8__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10066\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10126\,
datad => N_61587_I_0);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIMBLE_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_13__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10061\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10121\,
datad => N_61587_I_0);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_3_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000001")
port map (
combout => N_65775_RETI,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_13__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_11__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_5__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_9__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_17__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_15__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIGJKE_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_10__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10064\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10124\,
datad => N_61587_I_0);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIIO9M_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_2__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10072\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10132\,
datad => N_61587_I_0);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_COUNTSUCCESSIVEZERO36_SUB: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => N_65496_RETI,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_10__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_3__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_4__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_12__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_14__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_2__G2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_40_RNIBT6P1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000fcf0fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
dataf => N_65771_RETO,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_14_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(14),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_14__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(14));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNIRSLO_14_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fefcfaf0eeccaa00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349_RETI\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_DIVMULTV\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(14));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_35_RNITM313: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"abab0000ab000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO\,
dataa => CPI_D_INST_RETO(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_29_RNI6N313: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aabb0000a0b00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO\,
dataa => CPI_D_INST_RETO(12));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_22_RNI2OGP2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO\,
dataa => CPI_D_INST_RETO(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_16_RNIOPTH2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf000022230000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO\,
dataa => CPI_D_INST_RETO(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_RNIBJD01_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000004444404")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_3_RNIUG993: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f0000000d")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIOO9M_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_5__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10069\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10129\,
datad => N_61587_I_0);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIMO9M_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_4__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10070\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10130\,
datad => N_61587_I_0);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIKO9M_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_3__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10071\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10131\,
datad => N_61587_I_0);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M11S4: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7352_RETI\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_3__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_4__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_6__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_5__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(13),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_9_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(9),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(11),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_11__I0_I_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_1__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_16_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(10),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_16__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"faf0fefcaa00eecc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_RETI\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(375),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_142_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(142),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_14\(142),
datae => \GRLFPC2_0.FPO.FRAC\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNI8S1T_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"88088000ff7ff777")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10552\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10545\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10546\,
datac => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNI4HVV1_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0f000f00f0fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(45),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1\(45),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(19));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_42_RNIO38J_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5346\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_42_RNIO38J: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5346\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNII0D8_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ff000000ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNI1P63_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10545\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIT073_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10546\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_36_RNI41D81: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff8a800000757")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5410\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.EXTEND.TEMP_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIANGK_230_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcccf000cccc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.EXTEND.TEMP_0\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5346\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(230));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_36_RNIUQ6A1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffeca00000135f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5391\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.EXTEND.TEMP_0\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIIGIN1_186_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0ccaaaa0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1\(45),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(186));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNICDLR1_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"acac5353ff0000ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10746\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIITLR1_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"caca3535ff0000ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10744\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_48: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000780000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_48\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_20\,
datae => N_65707,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_16\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(35),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_63_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff2000ffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2\,
dataf => N_65610,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_2\,
datad => N_28250_2,
datac => N_28242,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_BUSYMULXFF_UN2_TEMP_SUB: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff75ffffff")
port map (
combout => N_65602,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3924\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3926\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.BUSYMULXFF.UN2_TEMP_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_O2_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff101010ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8573\,
dataf => N_32782_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9503\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9598\,
datac => N_34047_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0004")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_12\,
dataf => N_33652,
datae => N_33666,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_603\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff10000fff00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1027\,
dataf => N_33607_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9498\,
datad => N_33718_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9479\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff40000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_2\,
dataf => N_34330,
datae => N_32861_1,
datad => N_34341_1,
datac => N_32908_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffff80ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_7\,
dataf => N_32783,
datae => N_32844_2,
datad => N_32731,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_8_0\(47),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0400")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_9\,
dataf => N_32914,
datae => N_32907,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_26_1\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_4_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fff0fff07770fff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_4\(60),
dataf => N_33138_1,
datae => N_28921_1,
datad => N_33727_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A28_8_0\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff700070007000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_0\(8),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9522\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9523\,
datad => N_28312_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1734\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff404040ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9600\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1659\,
datad => N_33081_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff2000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_6\,
dataf => N_34181,
datae => N_34183,
datad => N_34263_2,
datac => N_28658_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffb000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_13\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_2\,
datad => N_32723_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_32_1\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f2002200f0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_0\,
dataf => N_33607_1,
datae => N_32859_1,
datad => N_32791_1,
datac => N_33984_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_44_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_44__G2_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9498\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9490\,
datad => N_32818_I,
datac => N_32974_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_4_2_RNIAP3P4_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff8000008080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_5\,
dataf => N_29653_1,
datae => N_32723_1,
datad => N_34059_1,
datac => N_34043_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_18_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffef000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_18\(60),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_2\(60),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_8\(60),
datad => N_34029,
datac => N_33738_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_11_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0d0f0d0f0ddfdd")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_11\(60),
dataf => N_29262_1,
datae => N_34341_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_1_TZ\(60),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A28_7_0\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_9\,
dataf => N_33902,
datae => N_33914,
datad => N_33735_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_10_0\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff40")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_7\,
dataf => N_33905,
datae => N_33899,
datad => N_33908,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11_1\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff4000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_10\,
dataf => N_33658,
datae => N_33653,
datad => N_33725_1,
datac => N_28652_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f2f02200f0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_13_0\,
dataf => N_33175,
datae => N_33222_2,
datad => N_33111,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A32_8_0\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_13_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00d00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_10\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_2\,
datae => N_33297_1,
datad => N_29366_1,
datac => N_28212_1_0,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff000f100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_17\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_10\,
datae => N_29262_1,
datad => N_33498_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A32_18_1\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_14_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A32_3_1\(57),
datae => N_32979_1,
datad => N_28227_1,
datac => N_32959_I,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_13_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbbbf000f000f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_5\,
dataf => N_33146_1,
datae => N_32789_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_A28_6_0\(56),
datac => N_33360_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_12_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000f000f222f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_11\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_603\,
datae => N_33725_1,
datad => N_33193,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_A28_5_1\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff40")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_10\,
dataf => N_33834,
datae => N_33827,
datad => N_33841,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_7_1\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff11001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_5\,
dataf => N_33503,
datae => N_32730_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_3_0\(52),
datac => N_33734_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff0004000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_11\,
dataf => N_33500,
datae => N_33727_2,
datad => N_28250_2,
datac => N_33899_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff8000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_15\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_10\,
datad => N_28212_1,
datac => N_33501_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0400")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_659\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1482\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9486\,
datac => N_29071_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_45_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff80")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9157\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9158\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9095_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_9_2_RNIBFN8D_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff1000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_2\,
datae => N_33291,
datad => N_33447_1,
datac => N_33293_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff8080ff80")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_9\,
dataf => N_33588,
datae => N_33193,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_27_0\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_23_0\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff4f0f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_6\,
dataf => N_33371,
datae => N_28921_1,
datad => N_28227_1,
datac => N_33365,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffff404040")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_974\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9523\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9517\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_1\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff10")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_6\,
dataf => N_32848,
datae => N_33079,
datad => N_33069,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_8_0\(18),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_5\,
dataf => N_33081,
datae => N_33068,
datad => N_33004,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_4_TZ\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_14_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffe000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_14__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9062\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_14__G2_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9502\,
datac => N_28222_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fdddf000f000f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9498\,
datae => N_28222_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1736\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_3_RNIR09D6_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff4000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_3\,
dataf => N_33783,
datae => N_33780,
datad => N_32786_1,
datac => N_33769,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_12_RNIS5QF6_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff00e0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_9\,
dataf => N_34056,
datae => N_34051,
datad => N_29653_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7_3_0\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff01000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_0\,
dataf => N_32842,
datae => N_29653_1,
datad => N_33368_1,
datac => N_32738_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff1000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_0\,
datad => N_28492_1,
datac => N_32831,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f010f00010100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_11\,
dataf => N_28212_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_6_1_0\(51),
datad => N_34343_1,
datac => N_33738_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83));
GRLFPC2_0_COMB_UN1_R_A_RS1_1_0_A2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"8808000000000000")
port map (
combout => \GRLFPC2_0.N_1841\,
dataf => \GRLFPC2_0.N_202\,
datae => \GRLFPC2_0.R.A.RS1D\,
datad => \GRLFPC2_0.R.STATE_O\(1),
datac => \GRLFPC2_0.R.STATE_O\(0),
datab => \GRLFPC2_0.COMB.FPDECODE.ST_O\,
dataa => N_155);
GRLFPC2_0_COMB_V_A_SEQERR_1_0_A2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000080000000000")
port map (
combout => \GRLFPC2_0.N_138\,
dataf => \GRLFPC2_0.N_90\,
datae => \GRLFPC2_0.FPCI_O\(59),
datad => \GRLFPC2_0.FPCI_O\(62),
datac => \GRLFPC2_0.FPCI_O\(69),
datab => \GRLFPC2_0.FPCI_O\(60),
dataa => \GRLFPC2_0.N_1837_O\);
\GRLFPC2_0_R_I_RES_RNO_63_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"5702ff005d08ff00")
port map (
combout => \GRLFPC2_0.COMB.V.I.RES_1\(63),
dataf => \GRLFPC2_0.FPI.OP2\(63),
datae => \GRLFPC2_0.N_1438_15\,
datad => \GRLFPC2_0.FPO.SIGN\,
datac => N_130,
datab => N_129,
dataa => N_13);
GRLFPC2_0_COMB_V_I_RDD_1_I_A3_15: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"8000000000000000")
port map (
combout => \GRLFPC2_0.N_1438_15\,
dataf => \GRLFPC2_0.COMB.V.I.RDD_1_I_A3_15_8\,
datae => \GRLFPC2_0.COMB.V.I.RDD_1_I_A3_15_9\,
datad => \GRLFPC2_0.COMB.V.E.FPOP_1\,
datac => \GRLFPC2_0.COMB.V.I.RDD_1_I_A3_15_7\,
datab => \GRLFPC2_0.FPCI_O\(62),
dataa => \GRLFPC2_0.FPCI_O\(60));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN12_SRTOSTICKY_1_RNIK26T: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"8888888888888880")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN12_SRTOSTICKY_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_4: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0087870000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTABORTNULLEXC_RNI04JG7: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0000000e0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_N_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_M2_E_RNIKOJ5843_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000f00f0f0fff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_N_6\,
dataf => D_N_7,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\,
datad => N_65488,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_2_RNI5G7A: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
dataf => N_65496,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_0\,
datac => N_65775);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA_SUB: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff00ffff0000")
port map (
combout => N_65549,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\,
datae => N_65719,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA_SUB_SUB: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff7f")
port map (
combout => N_65719,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_49_I\,
datae => \GRLFPC2_0.FPI.LDOP_0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_47: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000003c000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_47\,
dataf => N_65709,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_12\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_14\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_47_SUB: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fefbfdf7efbfdf7f")
port map (
combout => N_65709,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(28),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(14),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(14));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_48_SUB: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fefbefbffdf7df7f")
port map (
combout => N_65707,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(52),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(26),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(52));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_50_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3740088000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_42\,
dataf => N_65705,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_50_RNO_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f0f0000f0f000")
port map (
combout => N_65705,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(32));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_51_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3740088000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_44\,
dataf => N_65701,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(50),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_51_RNO_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f00f00f00f000")
port map (
combout => N_65701,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(42),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff0f0000fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10936\,
datae => N_65677,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_SUB_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000a500c300a500")
port map (
combout => N_65677,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN13_RESVEC\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(241));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_114_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0aaaae2aa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(114),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0_N_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0_M3_I_A3_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_115_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0aaaae2aa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(115),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0_N_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0_M3_I_A3_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(115));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_NOINSTANDNOEXC_0_A2_0_2_RNIFNJ9V: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff3f0ffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_51_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_877_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_551\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CONDMUXMULXFF_UN4_NOTSQRTLFTCC_I_O2_RNITCUV7: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff0f0f03cf0f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_663\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffdfffdfdfdff")
port map (
combout => N_65612,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datae => N_33507_1,
datad => N_33503_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffff0ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_0\,
datae => N_65612,
datad => N_33027,
datac => N_33031);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff85ffffffffffff")
port map (
combout => N_65611,
dataf => N_28549_1,
datae => N_28250_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff3")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_18\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_15\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_11\,
datad => N_33514,
datac => N_33504,
datab => N_65611);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_63_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000dfff")
port map (
combout => N_65610,
dataf => N_28254,
datae => N_28253,
datad => N_28243,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A14_0_S_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0f0ff0ffff")
port map (
combout => N_65608,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000f000")
port map (
combout => N_32838,
dataf => N_33004,
datae => N_65608,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81));
GRLFPC2_0_COMB_UN8_CCV_0_S: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000077707770777")
port map (
combout => N_65607,
dataf => \GRLFPC2_0.R.I.EXEC\,
datae => \GRLFPC2_0.R.I.INST\(19),
datad => \GRLFPC2_0.R.X.LD\,
datac => \GRLFPC2_0.R.X.AFSR\,
datab => \GRLFPC2_0.R.X.FPOP\,
dataa => N_348);
GRLFPC2_0_COMB_UN8_CCV_0_S_RNIHKLN: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000ccc0ccc0ccc")
port map (
combout => CPO_CCVZ,
dataf => N_279,
datae => \GRLFPC2_0.R.M.FPOP\,
datad => \GRLFPC2_0.R.E.FPOP\,
datac => N_210,
datab => N_65607);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_90_RNO_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f000f0f00000000")
port map (
combout => N_65588,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_A2_1_A2_9\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_A2_7_2\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1509\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIHHQ91_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000fff0fffffffff")
port map (
combout => N_65578,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(57));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_90_RNO_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cff0cff0cfffcff")
port map (
combout => N_65572,
dataf => \GRLFPC2_0.FPO.FRAC\(54),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_O2_0_RNIC6UT3_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcfffffff0f0f0f0")
port map (
combout => N_65570,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_TZ_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_402\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_551\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => N_59);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_M2_E_RNIKOJ5843: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000f00f0f0fff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1\,
dataf => D_N_7,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\,
datad => N_65488,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_83_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000fffff070")
port map (
combout => N_58999,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0_N_5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0_M3_I_A3_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0f0f0303030f03")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
dataf => N_27316,
datae => N_27258,
datad => N_27315,
datac => N_65549,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_2_IV_RNO_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f4f4f4f0f4")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_I_M\(12),
dataf => N_27316,
datae => N_27258,
datad => N_27315,
datac => N_65541,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN18_LOCOV_RNI2D3459: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0035ffffffffffff")
port map (
combout => N_65488,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_D\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0_0\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0\(9),
datac => N_27258,
datab => N_27310,
dataa => N_27309);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_53: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0080000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_53\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_40\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_24\,
datad => N_65528,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_4\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_6\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_7\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_53_SUB: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fefbefbffdf7df7f")
port map (
combout => N_65528,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(37),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(37));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_53_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"5720088000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_40\,
dataf => N_65526,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(43),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_53_RNO_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f00f00f00f000")
port map (
combout => N_65526,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(38),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff0f0000fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10934\,
datae => N_65522,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_SUB_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fa050000cc330000")
port map (
combout => N_65522,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fffa0000fefe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM12\,
datae => N_65516,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7778\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7777\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNII532TQ2_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fafaee445050ee44")
port map (
combout => N_53932,
dataf => N_27316,
datae => N_27258,
datad => N_27315,
datac => N_27314,
datab => N_27313,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN25_LOCOV_0_RNITQBF: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000004040000040c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0_0\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.REEXCOVUV.UN25_LOCOV_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(12),
datad => \GRLFPC2_0.FPO.EXP\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff30ffcfffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(27),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(30),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(28),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A8_2_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330cf00000000000")
port map (
combout => N_28252,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A8_2_0\(62),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_11_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3303303030000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_18_TZ\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_0_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f00000ff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_493\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_5\,
dataf => N_33353,
datae => N_29653_1,
datad => N_33055,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
GRLFPC2_0_R_I_EXEC_RNO_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000a800")
port map (
combout => \GRLFPC2_0.R.I.EXEC_0_0_G1_0_7945_I_3\,
dataf => \GRLFPC2_0.N_1438_15\,
datae => N_37320,
datad => N_37317,
datac => \GRLFPC2_0.R.X.FPOP\,
datab => \GRLFPC2_0.R.I.EXEC\,
dataa => N_11);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"08000800aaaa0800")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0_1\(37),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8524\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00aafcfc00aa0c0c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10085\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9789\,
datae => \GRLFPC2_0.FPI.LDOP_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(165),
dataa => N_703);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00aafcfc00aa0c0c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10101\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9805\,
datae => \GRLFPC2_0.FPI.LDOP_0_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(149),
dataa => N_719);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14_142_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300aaaafc00aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_14\(142),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(376),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(374),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(144));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccaaaaf0f0ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(25),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_15_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00aaaaccccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(15),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff000000ff484848")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_571\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9598\,
datad => N_33369_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_46_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0ccccaaaaff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(46),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaccccf0f0ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(50),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_17_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"1000000000000000")
port map (
combout => N_33845,
dataf => N_33734_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_1_A3_0_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fefe7efeffff7fff")
port map (
combout => N_28511,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1633\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_492\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_M2_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bfffffffbfff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_451\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_446\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(250),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(255),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(254),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(253),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_I_O2_4_4\(4));
GRLFPC2_0_COMB_LOCKGEN_UN8_DEPCHECK_RNI6D113: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0e0e00000f0e0f0e")
port map (
combout => \GRLFPC2_0.N_3477_1_I\,
dataf => \GRLFPC2_0.N_1714_I\,
datae => \GRLFPC2_0.N_1093\,
datad => \GRLFPC2_0.N_3458\,
datac => \GRLFPC2_0.N_1072\,
datab => \GRLFPC2_0.COMB.FPDECODE.ST\,
dataa => \GRLFPC2_0.N_951\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_23_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0aaaaccccff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(23),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_35_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0aaaaff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(35),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0aaaaff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(34),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00aaaaf0f0cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(39),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47));
\GRLFPC2_0_R_FSR_FTT_RNO_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000c480c4c0")
port map (
combout => \GRLFPC2_0.R.FSR.FTT_0_0_2__G1\,
dataf => \GRLFPC2_0.N_1015\,
datae => \GRLFPC2_0.N_58\,
datad => \GRLFPC2_0.R.X.SEQERR\,
datac => \GRLFPC2_0.R.FSR.FTT\(2),
datab => N_11,
dataa => \GRLFPC2_0.N_1105\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNI8IAN_247_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00807fffffffff")
port map (
combout => N_35132,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(247),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(249));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fdfdffccfdfd3300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fdfffdccfd33fd00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(52),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_44_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3bff08ff3b000800")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(44),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(44),
datae => N_53986,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_8_0_A2_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9498\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_3_0_A2_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9523\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_0_0_A2_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9600\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_8_2_0_A2_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9566\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_16_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1757\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_30_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1607\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_3_0_A2_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9598\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_17_1_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f00000000000")
port map (
combout => N_34272_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_1_1_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000c0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_1_1\(33),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_0_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0000000f000f00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_467\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_8_0_A2_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9511\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_1_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c0cc0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1200\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9486\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_0_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000c00000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0_0\(10),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_33_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1736\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_5_0_A2_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000f000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9502\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_0_A2_6: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000f00ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1758\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_13_0_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f0000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9492\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O23_0_0_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_0_0\(31),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_8_1_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f0000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_8_1\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O17_3_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c003c003f000000f")
port map (
combout => N_33276,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_4_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c0000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1049\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_467\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_3_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_661\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_15_I_O2_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ffffffffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_648\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_20_2_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000f")
port map (
combout => N_34047_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_2_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f00000f00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1713\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A21_0_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A21_0\(51),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_4_0_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000f0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A9_4_0\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A24_0_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A24_0\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_O28_8_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000f0000f0f0f")
port map (
combout => N_33710,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_10_2_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00000000000000")
port map (
combout => N_34335_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_14_3_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000f000000000")
port map (
combout => N_34339_3,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_14_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000030000")
port map (
combout => N_33842,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O8_2_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000f0000f000f0f")
port map (
combout => N_28242,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_0_2_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000ff")
port map (
combout => N_32722_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A32_8_0_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A32_8_0\(57),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_8_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000c00000000")
port map (
combout => N_34333,
dataf => N_32859_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_29_RNIB6P5A: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000f0ff000000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_5_TZ\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_0_1_0_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000c3f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0_1\(51),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_18_1_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000ff0000")
port map (
combout => N_34343_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_18_3_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff000000")
port map (
combout => N_32796_3,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_6_1_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f030c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_6_1\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_9_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000f0000000000")
port map (
combout => N_33795,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A32_18_1_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000c0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A32_18_1\(57),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_12_1_0_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_4_1\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A26_7_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3c0000000000000")
port map (
combout => N_33972,
dataf => N_34007,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A11_1_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fffc00000000000")
port map (
combout => N_28207,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A32_1_0\(57),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_10_TZ_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff3330fff0fff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_10_TZ\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_21_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => N_33229,
dataf => N_29653_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_10_2_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f000000000000")
port map (
combout => N_33838_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f000ffff00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_11_TZ\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff03ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_3\,
dataf => N_32792,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_2_0_0\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_5_1_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_A28_5_1\(56),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A28_4_1_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000003000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A28_4_1\(60),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A32_8_1_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000fff0")
port map (
combout => N_33222_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_4_2_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000ff00f0")
port map (
combout => N_34043_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A32_19_0_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000f00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A32_19_0\(57),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A11_5_3_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3f33000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A11_5_3\(61),
dataf => N_28211_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_O28_5_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff00ff")
port map (
combout => N_33193,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_1_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f00000ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_811\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_1_TZ_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0cffffff0cffcf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_1_TZ\(60),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_1_1_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff0000000000")
port map (
combout => N_34040_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_43_RNIGB99B: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000030300300333")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_13_TZ\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_5_0_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_16_0\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A14_2_2_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff000000")
port map (
combout => N_32840_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_7_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0c0000000c000c")
port map (
combout => N_28227,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A11_1_0_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A32_1_0\(57),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_12_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000030000")
port map (
combout => N_34051,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_16_0_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000f0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_32_1\(58),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_52_1_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_52_1\(58),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_4_0_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f000000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_4_0\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A32_28_2_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000ff0000")
port map (
combout => N_33152_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_O2_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff000000ff00ffff")
port map (
combout => N_33560,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A26_23_4_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000f0")
port map (
combout => N_33988_4,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_13_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000030000000")
port map (
combout => N_32735,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_42_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000003000")
port map (
combout => N_33444,
dataf => N_33111,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_0_0_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_0_0\(31),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_13_0_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_13_0\(51),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_11_2_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000f000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1592\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_2_1_RNIP800P_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff000f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_475\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_458\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_426\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_1_I_O2_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_812\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_12_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000300000000000")
port map (
combout => N_33220,
dataf => N_32818_I,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_7_3_0_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7_3_0\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_10_0_A2_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9509\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_13_0_A2_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000f00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9547\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_2_0_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_2_0\(31),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000c00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1133\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_467\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_3_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1031\,
dataf => N_32738_2,
datae => N_32738_1_0,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_32_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1734\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_35_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1749\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A2_8_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000ff")
port map (
combout => N_33756,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A11_2_2_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000f0000")
port map (
combout => N_28208_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_3_1_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03000000030f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_3_1\(32),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_11_0_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_11_0\(51),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A11_3_1_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A11_3_1\(61),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_12_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000000000")
port map (
combout => N_33175,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_2_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c00cc00000000")
port map (
combout => N_34041,
dataf => N_32738_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_6_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"300c000000000000")
port map (
combout => N_28226,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A28_7_0_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f00000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A28_7_0\(60),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_8_0_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f000f0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_8_0\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_2_0_A2_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9514\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_13_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000003000000000")
port map (
combout => N_34194,
dataf => N_29262_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_3_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000030000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9607\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_604\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_16_1_I_O2_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffff00ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_816\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O15_2_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff00ff00")
port map (
combout => N_33010,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_3_I_O2_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_814\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_1_A2_0_46_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000f00000f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1659\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_10_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000c00c0")
port map (
combout => N_32732,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_10_2_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff0000ff00")
port map (
combout => N_32732_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_9_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000030c000000000")
port map (
combout => N_32787,
dataf => N_33297_1,
datae => N_33004,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A11_5_2_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0000000f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A11_5_2\(61),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_18_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000c0000")
port map (
combout => N_33589,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_36_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c00000000000c0")
port map (
combout => N_33365,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000c00c00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1389\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A26_12_0\(11),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_13_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000c0000000000")
port map (
combout => N_34052,
dataf => N_28266_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_16_2_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff0000000000")
port map (
combout => N_34055_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_7_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000c00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_907\,
dataf => N_33340_I,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000ff0000")
port map (
combout => N_28263,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_10_I_O2_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff00ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_809\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_A2_34_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1672\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_3_0_A2_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000f00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9522\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_23_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000300000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1302\,
dataf => N_34029,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_9_I_O2_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0fffffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_525\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_14_2_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11810_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_0_0_A2_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9486\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_9_0_A2_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9517\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_1_35_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000030000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9200\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11641\,
datae => N_28266_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_14_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000030000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9373\,
dataf => N_28857_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_0\,
datad => N_32738_1_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A17_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000f0000000000")
port map (
combout => N_33283,
dataf => N_33278,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_4_1_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000ff0000")
port map (
combout => N_28312_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_0_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000003000003000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffcfff30ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(19),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(37),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff30ffcfffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(56),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_20_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffcfff30ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(20),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(36),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(37),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_21_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffcfff30ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(21),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(35),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_22_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff30ffcfffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(22),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(35),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_23_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffcfff30ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(23),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(33),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffcfff30ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(24),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffcfff30ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(26),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(30),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffcfff30ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(54),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff30ffcfffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(36),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(21),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffcfff30ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(53),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffcfff30ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(9),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(10),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffcfff30ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(52),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffcfff30ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(51),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffcfff30ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(50),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffcfff30ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(49),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(50),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff30ffcfffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(8),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(49),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_22_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0ff0f000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(22),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(22),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(21),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
GRLFPC2_0_R_A_FPOP_RNIE2QG: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
combout => \GRLFPC2_0.COMB.V.E.FPOP_1\,
dataf => \GRLFPC2_0.R.A.FPOP\,
datae => N_156,
datad => N_157);
GRLFPC2_0_R_E_LD_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
combout => \GRLFPC2_0.R.E.LD_0_0_G1\,
dataf => \GRLFPC2_0.R.A.LD\,
datae => N_156,
datad => N_157);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_10_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000c000000")
port map (
combout => N_32788,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_1_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10859\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_1_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff000000fff00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10860\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_1_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10864\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_1_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10862\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_13_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000c000000000")
port map (
combout => N_33841,
dataf => N_28549_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_5_1_0_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000c0000003f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_5_1\(59),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_6_1_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f000f000f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_6_1\(59),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_20_1_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f00000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_4_1\(59),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_6_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3f00000000000000")
port map (
combout => N_32976,
dataf => N_32861_1,
datae => N_32738_2,
datad => N_32738_1_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_26_1_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c0c0c00000c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_26_1\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_3_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccfff000cc00f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(238),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(251));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_5_0_A2_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9503\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A28_0_1_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000c0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A28_0_1\(60),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_5_0_A2_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9525\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_O23_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff000000ffff00ff")
port map (
combout => N_33870,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_20_1_I_O2_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fffffffffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_571\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_3_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1236\,
dataf => N_28266_2,
datae => N_32738_1_0,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_7_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c0000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1206\,
dataf => N_33070_1,
datae => N_28266_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_8_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1036\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11641\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\,
datad => N_34263_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_17_1_0_A2_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9479\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cc000000fc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW_6\(0),
dataf => N_61,
datae => N_65,
datad => N_64,
datac => N_60,
datab => N_62);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f00000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7260\,
dataf => N_60,
datae => N_65,
datad => N_62,
datac => N_64);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7259\,
dataf => N_60,
datae => N_65,
datad => N_62,
datac => N_64);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_1_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0f0000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10857\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_1_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10858\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_33_0_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000f0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_33_0\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_25_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000330f0000")
port map (
combout => N_33427,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_782\,
datae => N_32727_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_M2_0_O2_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8619\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIGNP91_247_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffc00000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_893\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1637\,
datae => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(247),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(249));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_0_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333cccc0ff00ff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CHECKOVANDDENORM_UN13_NOTPOSSIBLEOV_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff000000c0c0c0c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_0\,
dataf => N_27258,
datae => N_27302,
datad => N_27298,
datac => N_27301,
datab => N_27297);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CHECKOVANDDENORM_UN13_NOTPOSSIBLEOV_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f00000cc00cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_1\,
dataf => N_27258,
datae => N_27304,
datad => N_27303,
datac => N_27296,
datab => N_27295);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_24: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"003f3f0000c0c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_24\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(46),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_41_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => N_33658,
dataf => N_32861_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A28_16_3_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000f000000000")
port map (
combout => N_33735_3,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_4_0_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c3c3c3c00ffff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_20: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03ff30000c00c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_20\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_15_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000300000000000")
port map (
combout => N_33514,
dataf => N_29262_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_11_1_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000030030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11_1\(59),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_27_0_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f0000030f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_27_0\(27),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_1_1_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000ff")
port map (
combout => N_34256_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_4_2_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000f00000")
port map (
combout => N_32974_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_16_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000003000000000")
port map (
combout => N_32794,
dataf => N_32730_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O2_0_0_A2_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1595\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_7_A2_0_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f0000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1586\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_1_0_A2_44_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000030000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9095_1\,
dataf => N_34263_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_40_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000000000")
port map (
combout => N_33369,
dataf => N_33984_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_7_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000030000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8834\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datae => N_34263_2,
datad => N_28266_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_2_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9645\,
dataf => N_33070_1,
datae => N_34263_2,
datad => N_32818_I,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_40_1_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => N_33369_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_18_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1714\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_20_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1800\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_28: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"003f3f0000c0c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_28\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(39),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(30),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A8_2_0_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A8_2_0\(62),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff9f0f9b00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_15\,
dataf => N_32797,
datae => N_33718_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_1_1\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_36_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3fff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1493\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_875\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_44_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000c00000000000")
port map (
combout => N_33661,
dataf => N_28250_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_28_1_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f00ff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_28_1\(58),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_8_0_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000f0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_8_0\(18),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_7_0_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7_0\(52),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A23_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fccc00000000")
port map (
combout => N_33498,
dataf => N_33498_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_604\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_3_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33000000000000")
port map (
combout => N_33899,
dataf => N_33659_1,
datae => N_33899_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_15_2_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000000000000000")
port map (
combout => N_34340_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_2_1_0_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33000f0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_2_1\(59),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A32_15_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00003c0000000000")
port map (
combout => N_33139,
dataf => N_28271_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_603\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_604\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83));
\GRLFPC2_0_R_STATE_RNIVPL21_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcfffffffcfffc")
port map (
combout => \GRLFPC2_0.N_67\,
dataf => \GRLFPC2_0.R.STATE\(0),
datae => \GRLFPC2_0.R.STATE\(1),
datad => N_88,
datac => N_14,
datab => N_87);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_7_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000c")
port map (
combout => N_33578,
dataf => N_33984_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_12_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000000000")
port map (
combout => N_34337,
dataf => N_33436_1,
datae => N_32859_1,
datad => N_28251_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_16_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000c000000000")
port map (
combout => N_34271,
dataf => N_33070_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_19_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0003000000000000")
port map (
combout => N_33518,
dataf => N_33070_1,
datae => N_33984_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A26_1_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000ff")
port map (
combout => N_34133_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_16_2_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000f000")
port map (
combout => N_33718_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A26_17_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000c0000000000")
port map (
combout => N_33982,
dataf => N_33734_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A26_3_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000003000000")
port map (
combout => N_33968,
dataf => N_33074_1,
datae => N_34263_2,
datad => N_33179,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_14_S_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f000000030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_A2_14_S\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1566\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1618\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(66));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A26_5_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333c000000000000")
port map (
combout => N_33970,
dataf => N_33507_1,
datae => N_28251_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN3_INEXACT: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000030033")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4664\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_28: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0003000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_28\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_26\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_20\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_43_1_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9490\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_37_1_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f00000000")
port map (
combout => N_33373_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_11_0_O2_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffff0ffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_473\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1194\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_2_1_RNIBS5F9_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f303f00003030000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_426\,
dataf => N_32782_1,
datae => N_33725_1,
datad => N_34329_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_20_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000003000000")
port map (
combout => N_33916,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11641\,
datae => N_29195_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A2_8_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000ff0000")
port map (
combout => N_33253,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_14_1_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000f0")
port map (
combout => N_34059_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_23_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1301\,
dataf => N_32844_2,
datae => N_33070_1,
datad => N_34263_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_1_23_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000300000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1303\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_782\,
datae => N_32738_1_0,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_4_1_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000c0000c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_4_1\(33),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_1_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000c000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1135\,
dataf => N_32844_2,
datae => N_33070_1,
datad => N_34263_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_5_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1191\,
dataf => N_34263_2,
datae => N_32738_1_0,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_2_30_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1222_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_20_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000c0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1304\,
dataf => N_33074_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_797\,
datad => N_33263_I,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_9_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000c00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1054\,
dataf => N_33074_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_9_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9418\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\,
datad => N_33607_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_24_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8941\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_4_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000c0000000000")
port map (
combout => N_32974,
dataf => N_32844_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11641\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_0_1_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f00000f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_0_1\(13),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_15_2_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ff00")
port map (
combout => N_28390_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_2_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000c")
port map (
combout => N_34327,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_797\,
datae => N_34311_I,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_19_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1482\,
dataf => N_33074_1,
datae => N_32782_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_4_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000c000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1832\,
dataf => N_32782_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_4_37_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000c000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1588\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11641\,
datae => N_33074_1,
datad => N_32782_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_4_0_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_4_0\(12),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_6_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000c000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1697\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datae => N_33074_1,
datad => N_32782_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_X2_2_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0000000ff0f0f0")
port map (
combout => N_32956_I,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_11_0_A2_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c0000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9349\,
dataf => N_32844_2,
datae => N_32782_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_7_0_A2_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9099\,
dataf => N_32844_2,
datae => N_32782_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_A2_25_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000c00000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1768\,
dataf => N_32782_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_1_A2_41_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000c000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9165\,
dataf => N_33340_I,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_14_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => N_33081,
dataf => N_29262_1,
datae => N_33507_1,
datad => N_33004,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A28_8_2_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000ff0000")
port map (
combout => N_33727_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_6_1_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000003c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_6_1\(31),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_0_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f000f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_SA_I_1_0_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff3c3c00003c3c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1_0_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(316),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(258));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_1_RNI4IGM: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0f0c0c0c0c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1274_I\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10626\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(316));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_30_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000300000000000")
port map (
combout => N_33359,
dataf => N_32844_2,
datae => N_29195_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_12_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000003000")
port map (
combout => N_34123,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datae => N_32858_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_0_1_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => N_34325_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_38_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000300")
port map (
combout => N_32916,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11641\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_21_1_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => N_34132_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_1_0_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000030003000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_1\(26),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_9_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000c0")
port map (
combout => N_33683,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_10_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000c000000")
port map (
combout => N_34191,
dataf => N_33548,
datae => N_33340_I,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_13_1_0_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_13_1\(51),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_1_2_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ff00")
port map (
combout => N_34326_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIA1PQ_77_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffcccf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CONDMUXMULXFF_UN4_NOTSQRTLFTCC_I_O2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff0f0f0ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_663\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_0_A2_8_A0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f0f0f0ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1809\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_0_O2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0c0c0c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_551\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_479\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(63));
GRLFPC2_0_R_A_LD_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000c00")
port map (
combout => \GRLFPC2_0.R.A.LD_0_0_G1\,
dataf => \GRLFPC2_0.N_3477_1_I\,
datae => \GRLFPC2_0.N_67\,
datad => \GRLFPC2_0.R.A.LD_0_0_G1_3\,
datac => N_76,
datab => N_77);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_14_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f0f0fff0f0f0f")
port map (
combout => N_53873,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_16_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0f0f0f000f0f0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SCTRL_NEW\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNICR8O9O3_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff00fcfcfcfc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0\(9),
dataf => N_27258,
datae => N_27314,
datad => N_27312,
datac => N_27313,
datab => N_27311);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_31_RNIH52J_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000300030003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_389\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1677\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1770\,
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_O2_29_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffff0ffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_743\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
datae => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A11_3_0_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0000000f000f00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A11_3_0\(61),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_14_1_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0ff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_15_0\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNI9BPM_247_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000300000003fffc")
port map (
combout => N_35133,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(249),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(247));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_39_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => N_32917,
dataf => N_33447_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_44_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000003000000")
port map (
combout => N_33373,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datae => N_33607_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_4_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000c00")
port map (
combout => N_33071,
dataf => N_33146_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_604\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_42_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000c0000000000")
port map (
combout => N_33371,
dataf => N_33074_1,
datae => N_33548,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_0_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9369\,
dataf => N_33146_1,
datae => N_33798_I,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A2_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ff00")
port map (
combout => N_32789_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_32_1_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000c030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_32_1\(27),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_6_0_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000330f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_0_A28_6_0\(56),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_1_37_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0c0000cc000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0_1\(37),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_1_0_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_1_0\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_34_0_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000030000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_34_0\(58),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_11_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000300")
port map (
combout => N_32981,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_603\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A20_1_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000ff0000")
port map (
combout => N_32981_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A14_6_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000300000000000")
port map (
combout => N_32844,
dataf => N_32844_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_0\,
datad => N_32821,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_9_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000303300000000")
port map (
combout => N_32731,
dataf => N_32731_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_9_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000003000")
port map (
combout => N_33905,
dataf => N_33659_1,
datae => N_33004,
datad => N_28211_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_0_A28_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030cc0000000000")
port map (
combout => N_33207,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A32_19_0\(57),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_10_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000c0000000")
port map (
combout => N_34121,
dataf => N_28264_1,
datae => N_28730_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_17_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000030000000")
port map (
combout => N_34056,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_782\,
datae => N_32782_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_0_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f3330000")
port map (
combout => N_34111,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_719\,
datae => N_33447_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_33_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000030000000")
port map (
combout => N_33650,
dataf => N_32982_1,
datae => N_28492_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A28_19_1_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => N_33738_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_14_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => N_32792,
dataf => N_28658_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_46_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_46__G2\,
dataf => N_34029,
datae => N_33340_I,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_9_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000c00000")
port map (
combout => N_33076,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\,
datae => N_29262_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_13_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000c0000")
port map (
combout => N_33584,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_28_0_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff000f0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_28_0\(58),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_36_0_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_15_1\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14_172_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000003000000fc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_14\(172),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(376),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(374));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_T_3_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33333cfc33333c0c")
port map (
combout => N_53995,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(374),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(376),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(375),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(377));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_15_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000003000000")
port map (
combout => N_33911,
dataf => N_33004,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_16_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3033000000000000")
port map (
combout => N_33224,
dataf => N_33725_1,
datae => N_32909_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A11_4_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000300000000000")
port map (
combout => N_28210,
dataf => N_32844_3,
datae => N_32909_1,
datad => N_29195_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_36_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03000c0000000000")
port map (
combout => N_33653,
dataf => N_33503_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000b900")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_6\,
dataf => N_32727,
datae => N_33178,
datad => N_28261_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
GRLFPC2_0_COMB_FPDECODE_RDD5_0_A2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => \GRLFPC2_0.N_925\,
dataf => \GRLFPC2_0.N_3468\,
datae => N_59,
datad => N_58,
datac => N_63,
datab => N_64);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_8_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f0000000000000")
port map (
combout => N_33794,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_17_1_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff0000000000")
port map (
combout => N_33668_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_8_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000300000")
port map (
combout => N_34119,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_782\,
datae => N_29366_1,
datad => N_33734_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_52_0_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_52_0\(58),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000003000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9327\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_531\,
datae => N_33607_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_9_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => N_34120,
dataf => N_34029,
datae => N_28730_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_1_0_A2_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000300000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9397\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datae => N_33074_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_6_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000003000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_974\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_4_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000003000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1237\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11641\,
datae => N_33607_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_0_A2_7: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cf000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1769\,
dataf => N_33607_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(66),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(67));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_7_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1374\,
dataf => N_32844_2,
datae => N_32738_1_0,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_7_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1682\,
dataf => N_32844_2,
datae => N_33436_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_7_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000030000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9166\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11641\,
datae => N_33074_1,
datad => N_32782_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_3_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1648\,
dataf => N_33070_1,
datae => N_33074_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_2_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000300030000000")
port map (
combout => N_33830,
dataf => N_29653_1,
datae => N_33070_1,
datad => N_29518_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_34_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c0f0000000000000")
port map (
combout => N_32912,
dataf => N_33368_1,
datae => N_32727_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_35_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cf00000000000000")
port map (
combout => N_33652,
dataf => N_33652_1,
datae => N_33507_1,
datad => N_32909_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_14_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000300000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_948\,
dataf => N_33070_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_21_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => N_32946,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_30_RNIDO6R4_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff3000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_9\,
dataf => N_33432,
datae => N_33445,
datad => N_28857_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_2_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"030c000000000000")
port map (
combout => N_32972,
dataf => N_32844_3,
datae => N_32727_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A32_13_1_0_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000ffff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A32_13_1_0\(57),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
GRLFPC2_0_RS1D_CNST_0_A2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000c00000000000")
port map (
combout => \GRLFPC2_0.RS1D_CNST\,
dataf => N_84,
datae => N_75,
datad => \GRLFPC2_0.N_2888\,
datac => N_77,
datab => N_74);
GRLFPC2_0_RS1V12_TZ: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f00000000000f000")
port map (
combout => \GRLFPC2_0.RS1V12_TZ\,
dataf => N_72,
datae => N_73,
datad => N_77,
datac => N_74);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_16_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0003000000000000")
port map (
combout => N_33844,
dataf => N_33984_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_43_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => N_32921,
dataf => N_34329_1,
datae => N_33607_1,
datad => N_32796_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_19_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000000000")
port map (
combout => N_32797,
dataf => N_32730_1,
datae => N_32738_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_11_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000303300000000")
port map (
combout => N_33839,
dataf => N_33543,
datae => N_33178,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_4_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000030000300")
port map (
combout => N_33832,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_531\,
datae => N_32722_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_26_2_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
combout => N_32904_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A32_11_0_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000f00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A32_11_0\(57),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_3_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0c0c0000000000")
port map (
combout => N_33574,
dataf => N_28264_1,
datae => N_33146_1,
datad => N_29366_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A32_10_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f030000")
port map (
combout => N_33134,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_603\,
datae => N_28730_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_15_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0c000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_2\,
dataf => N_33149,
datae => N_33146_1,
datad => N_28250_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_31_RNI334M4_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0c000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_3\,
dataf => N_33433,
datae => N_33138_1,
datad => N_33146_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_20_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000000000")
port map (
combout => N_34059,
dataf => N_32782_1,
datae => N_28492_1,
datad => N_32738_1_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_5\,
dataf => N_33911,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_7_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000030000")
port map (
combout => N_32729,
dataf => N_33548,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_603\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_12_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000c")
port map (
combout => N_33079,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_603\,
datae => N_33004,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_13_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000030000")
port map (
combout => N_33297,
dataf => N_33548,
datae => N_33297_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_6_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030000000000000")
port map (
combout => N_33073,
dataf => N_28492_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_20_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000030000000000")
port map (
combout => N_32798,
dataf => N_33507_1,
datae => N_33004,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_7_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000000000")
port map (
combout => N_32785,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datae => N_33297_1,
datad => N_33734_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_38_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0c000000000000")
port map (
combout => N_33440,
dataf => N_33574_1,
datae => N_28658_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_45_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000000000")
port map (
combout => N_33447,
dataf => N_33574_1,
datae => N_33146_1,
datad => N_33447_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_31_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000003000000000")
port map (
combout => N_33648,
dataf => N_33735_1,
datae => N_32959_I,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_38_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000300000")
port map (
combout => N_33655,
dataf => N_33735_1,
datae => N_33734_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81));
\GRLFPC2_0_R_A_AFQ_RET_RNISCAR_9_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000f0f000000000")
port map (
combout => \GRLFPC2_0.R.E.AFQ_RET_0_0_G1_5\,
dataf => \GRLFPC2_0.FPCI_O\(69),
datae => \GRLFPC2_0.R.STATE_O\(0),
datad => \GRLFPC2_0.R.STATE_O\(1),
datac => \GRLFPC2_0.FPCI_O\(70));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A14_3_1_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c0cccc00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_3_1\(25),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_3_0_A2_44_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9157\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
datad => N_28857_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_8_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1053\,
dataf => N_33074_1,
datae => N_32782_1,
datad => N_32738_1_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_4_0_A2_44_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000c00000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9158\,
dataf => N_32844_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11641\,
datad => N_32782_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_40_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1278\,
dataf => N_32844_2,
datae => N_28266_2,
datad => N_32738_1_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_22_0_A2_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000c0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9062\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datae => N_28857_1,
datad => N_28266_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_5_44_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9159\,
dataf => N_33070_1,
datae => N_33074_1,
datad => N_32782_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A14_10_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => N_32848,
dataf => N_29653_1,
datae => N_33146_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_43_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => N_33445,
dataf => N_33081_1,
datae => N_28227_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_6_0_A2_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9570\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
GRLFPC2_0_R_E_SEQERR_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaa080000000000")
port map (
combout => \GRLFPC2_0.R.E.SEQERR_0_0_G1\,
dataf => \GRLFPC2_0.N_552_1_0\,
datae => \GRLFPC2_0.N_138\,
datad => \GRLFPC2_0.N_94\,
datac => \GRLFPC2_0.FPCI_O\(62),
datab => \GRLFPC2_0.FPCI_O\(69),
dataa => \GRLFPC2_0.FPCI_O\(70));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_9_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030000000000000")
port map (
combout => N_34334,
dataf => N_33543,
datae => N_29366_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_8_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => N_33904,
dataf => N_33140_1,
datae => N_33004,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A26_20_2_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000f")
port map (
combout => N_33985_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_14_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc00000000000000")
port map (
combout => N_33513,
dataf => N_29653_1,
datae => N_33725_1,
datad => N_33146_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_14_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0003000000000000")
port map (
combout => N_34195,
dataf => N_33659_1,
datae => N_28658_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_14_1_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000ff")
port map (
combout => N_34195_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A26_10_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0003000000000000")
port map (
combout => N_33975,
dataf => N_28211_1,
datae => N_34311_I,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A26_11_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000000000")
port map (
combout => N_33976,
dataf => N_32979_1,
datae => N_34311_I,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A28_8_0_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000f00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A28_8_0\(60),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN50_ZERO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33fffffffff0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6961\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN48_ZERO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33ffffffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN54_ZERO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000f33")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIN0DJ_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0ccf0ccf0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_372__G1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_16_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => N_34127,
dataf => N_33735_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_531\,
datad => N_32909_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A32_0_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c000000c0c00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A32_0\(57),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_18_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => N_33914,
dataf => N_33574_1,
datae => N_32727_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_17_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000c000")
port map (
combout => N_33225,
dataf => N_33055,
datae => N_33503_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_31_1_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => N_33360_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_34_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030000000000000")
port map (
combout => N_33363,
dataf => N_33055,
datae => N_28857_1,
datad => N_32821,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A28_10_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000300000000000")
port map (
combout => N_33729,
dataf => N_28634_1,
datae => N_33138_1,
datad => N_33503_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_O28_9_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff00ff00")
port map (
combout => N_33715,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff30000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_4\,
dataf => N_33139,
datae => N_33659_1,
datad => N_32909_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_10_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000030000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_8\,
dataf => N_33659_1,
datae => N_34341_1,
datad => N_28261_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A32_24_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000030000000")
port map (
combout => N_33148,
dataf => N_33548,
datae => N_29262_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIPHE9_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0fff0fff03f30")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0_M3_I_A3_0\,
dataf => \GRLFPC2_0.FPI.LDOP_1_2\,
datae => \GRLFPC2_0.R.MK.RST2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datab => N_11);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_64_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff33f3ffff3333")
port map (
combout => \GRLFPC2_0.FPI.RST\,
dataf => \GRLFPC2_0.R.MK.RST_4\,
datae => \GRLFPC2_0.R.MK.RST2\,
datad => \GRLFPC2_0.R.MK.RST2_O\,
datac => \GRLFPC2_0.COMB.ANNULFPU_1_O\,
datab => N_11);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN1_U_SNNOTDB: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00f0ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462\,
dataf => \GRLFPC2_0.FPI.LDOP_1_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.R.MK.RST2\,
datac => N_11);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNITSA8_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
dataf => \GRLFPC2_0.FPI.LDOP_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datad => \GRLFPC2_0.R.MK.RST2\,
datac => N_11);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNISSA8_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0fff")
port map (
combout => N_61587_I,
dataf => \GRLFPC2_0.FPI.LDOP_1\,
datae => \GRLFPC2_0.R.MK.RST2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(5),
datac => N_11);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIGEPD_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000f000")
port map (
combout => N_37019_2,
dataf => \GRLFPC2_0.FPI.LDOP_1\,
datae => \GRLFPC2_0.R.MK.RST2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datac => N_11);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_68_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\,
dataf => \GRLFPC2_0.FPI.LDOP_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(12),
datad => \GRLFPC2_0.R.MK.RST2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(47),
datab => N_11);
GRLFPC2_0_FPI_LDOP: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff00ff")
port map (
combout => \GRLFPC2_0.FPI.LDOP\,
dataf => \GRLFPC2_0.FPI.LDOP_1_2\,
datae => \GRLFPC2_0.R.MK.RST2\,
datad => N_11);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_4_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000300000000000")
port map (
combout => N_33900,
dataf => N_32859_1,
datae => N_33577_1,
datad => N_33734_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_16_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => N_33912,
dataf => N_33735_1,
datae => N_28921_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_10_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030000000000000")
port map (
combout => N_34049,
dataf => N_29653_1,
datae => N_32782_1,
datad => N_33899_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_6_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000003000000")
port map (
combout => N_34117,
dataf => N_34311_I,
datae => N_29518_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_0_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc33cc0f0ff0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A11_6_1_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ff00")
port map (
combout => N_28212_1_0,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_3_0_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_3_0\(51),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84));
GRLFPC2_0_COMB_ANNULFPU_1_U_0_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcfcfcff000000")
port map (
combout => \GRLFPC2_0.COMB.ANNULFPU_1_U_0_0\,
dataf => \GRLFPC2_0.R.E.FPOP\,
datae => \GRLFPC2_0.R.A.FPOP\,
datad => \GRLFPC2_0.N_1685\,
datac => N_225,
datab => N_226);
GRLFPC2_0_R_M_FPOP_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
combout => \GRLFPC2_0.R.M.FPOP_0_0_G1\,
dataf => \GRLFPC2_0.R.E.FPOP\,
datae => N_225,
datad => N_226);
GRLFPC2_0_R_M_LD_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
combout => \GRLFPC2_0.R.M.LD_0_0_G1\,
dataf => \GRLFPC2_0.R.E.LD\,
datae => N_225,
datad => N_226);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_5_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000003fffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_5\(60),
dataf => N_33733,
datae => N_33543,
datad => N_32859_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_7_37_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1718\,
dataf => N_33735_1,
datae => N_33074_1,
datad => N_34329_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_10_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1055\,
dataf => N_33735_1,
datae => N_33074_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_1_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c0000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1212\,
dataf => N_32844_2,
datae => N_34263_2,
datad => N_33652_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_2_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3f00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9371\,
dataf => N_33074_1,
datae => N_34263_2,
datad => N_33574_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33c0c00000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_5\,
dataf => N_32861_1,
datae => N_32982_1,
datad => N_33899_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00c00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_693\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8537\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8524\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_7_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000c0000000000")
port map (
combout => N_33903,
dataf => N_29195_1,
datae => N_33721_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_13_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => N_34268,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0300fcf0000")
port map (
combout => N_53985,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(56),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
GRLFPC2_0_R_A_FPOP_RNIUNSG: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.N_1714_I\,
dataf => \GRLFPC2_0.R.X.FPOP\,
datae => \GRLFPC2_0.R.I.EXEC\,
datad => \GRLFPC2_0.R.M.FPOP\,
datac => \GRLFPC2_0.R.E.FPOP\,
datab => \GRLFPC2_0.R.A.FPOP\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_0_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc33cc0f0ff0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_2_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c300000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1235\,
dataf => N_32844_2,
datae => N_34263_2,
datad => N_32796_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c300000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1744\,
dataf => N_32844_2,
datae => N_34341_1,
datad => N_32796_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_6_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9375\,
dataf => N_33074_1,
datae => N_34341_1,
datad => N_32796_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_9_2_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000ff0000")
port map (
combout => N_33293_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_4_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3003000000000000")
port map (
combout => N_34329,
dataf => N_29653_1,
datae => N_34329_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_30_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c00000000c0000")
port map (
combout => N_32908,
dataf => N_32844_2,
datae => N_28271_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A32_1_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ff00")
port map (
combout => N_33123_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_11_0_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f00000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_11_0\(32),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O17_4_RNIQ7IB5_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0c000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_4\,
dataf => N_33286,
datae => N_33277,
datad => N_33899_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_9_0_0_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000c000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_9_0_0\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN20_ZERO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fffffffffccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5771\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNI8KVE_23_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fffff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5452\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN18_ZERO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fffffffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN24_ZERO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000330f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23));
GRLFPC2_0_R_X_FPOP_RNINRLL: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0003000000000000")
port map (
combout => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
dataf => \GRLFPC2_0.R.X.FPOP\,
datae => N_13,
datad => N_364,
datac => N_363,
datab => N_14);
GRLFPC2_0_R_I_EXEC_RNO_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffc0000ffff0003")
port map (
combout => N_37317,
dataf => \GRLFPC2_0.R.X.SEQERR\,
datae => \GRLFPC2_0.R.I.EXEC\,
datad => N_364,
datac => N_363,
datab => N_14);
GRLFPC2_0_R_X_FPOP_RNIAQIJ: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f00000000")
port map (
combout => N_37343_I_0,
dataf => \GRLFPC2_0.R.X.FPOP\,
datae => N_364,
datad => N_363,
datac => N_14);
GRLFPC2_0_R_X_AFSR_RNI0Q3P: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0003000000000000")
port map (
combout => \GRLFPC2_0.N_1171\,
dataf => \GRLFPC2_0.R.X.LD\,
datae => \GRLFPC2_0.R.X.AFSR\,
datad => N_364,
datac => N_363,
datab => N_14);
GRLFPC2_0_WRADDR_0_SQMUXA: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000030000")
port map (
combout => \GRLFPC2_0.N_1243\,
dataf => \GRLFPC2_0.R.X.AFSR\,
datae => \GRLFPC2_0.R.X.LD\,
datad => N_364,
datac => N_363,
datab => N_14);
GRLFPC2_0_RS2_0_SQMUXA_0_0_A2_0_RNI8D6T: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000c000000")
port map (
combout => \GRLFPC2_0.N_3458\,
dataf => N_76,
datae => \GRLFPC2_0.N_45\,
datad => \GRLFPC2_0.N_3462\,
datac => N_74,
datab => N_83);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000c3000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1134\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11641\,
datae => N_33074_1,
datad => N_33734_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_24_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c3c3c30000000000")
port map (
combout => N_33353,
dataf => N_32738_1,
datae => N_32723_1,
datad => N_28921_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_2_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c300000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1201\,
dataf => N_32844_2,
datae => N_32738_1_0,
datad => N_33984_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
\GRLFPC2_0_COMB_RF1REN_1_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0fff0ffffff0000")
port map (
combout => RFI1_REN2Z,
dataf => N_398,
datae => \GRLFPC2_0.N_3150\,
datad => N_399,
datac => N_400);
GRLFPC2_0_WRADDR_0_SQMUXA_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
dataf => N_398,
datae => N_399,
datad => N_400);
GRLFPC2_0_COMB_V_FSR_RD_1_SN_M2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fffffff00000000")
port map (
combout => \GRLFPC2_0.N_3027\,
dataf => N_11,
datae => N_400,
datad => N_399,
datac => N_398);
GRLFPC2_0_V_FSR_CEXC_0_SQMUXA: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fffffff00000000")
port map (
combout => \GRLFPC2_0.V.FSR.CEXC_0_SQMUXA\,
dataf => \GRLFPC2_0.N_1439\,
datae => N_400,
datad => N_399,
datac => N_398);
GRLFPC2_0_V_STATE_1_SQMUXA: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3fff0000ffff0000")
port map (
combout => \GRLFPC2_0.N_1667\,
dataf => N_434,
datae => N_11,
datad => N_400,
datac => N_399,
datab => N_398);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_3_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c3000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1214\,
dataf => N_33070_1,
datae => N_32723_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_1_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff000000c3000000")
port map (
combout => N_33572,
dataf => N_28264_1,
datae => N_29071_1,
datad => N_28564_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN35_ZERO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33fffffffff0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6583\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f330000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5458\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN33_ZERO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33ffffffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN39_ZERO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000f33")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0300fcf0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(5),
dataf => N_53884,
datae => N_53883,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0300fcf0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(6),
dataf => N_53905,
datae => N_53925,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0300fcf0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(7),
dataf => N_53924,
datae => N_53926,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_9_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0fcff0300000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(9),
dataf => N_53929,
datae => N_53883,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(372));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIG40F_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f330000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5446\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN40_SHDVAR: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffe00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN40_SHDVAR\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5416\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_1_RNIO2GH: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f033ff330fcc00cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_12231\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(258));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_6_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000003000000000")
port map (
combout => N_33902,
dataf => N_33659_1,
datae => N_29366_1,
datad => N_32738_1_0,
datac => N_33734_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_14_RNI4K633_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00300000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_948\,
datae => N_33074_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\,
datac => N_34329_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_3_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000003c3f")
port map (
combout => N_34042,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_782\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c0000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1388\,
dataf => N_32844_2,
datae => N_28266_2,
datad => N_28251_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fccf00f33f0cc")
port map (
combout => N_53044,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c3f03cff3c0fc30")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0330f33ffccf0cc0")
port map (
combout => N_53175,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30cf03fc3fc0f30c")
port map (
combout => N_53198,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03fc30cff30c3fc0")
port map (
combout => N_53221,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30cf03fc3fc0f30c")
port map (
combout => N_53244,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0fc33c3cc3f0f0")
port map (
combout => N_53267,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0fc33c3cc3f0f0")
port map (
combout => N_53290,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0fc33c3cc3f0f0")
port map (
combout => N_53313,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0fc33c3cc3f0f0")
port map (
combout => N_53336,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0fc33c3cc3f0f0")
port map (
combout => N_52670,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0fc33c3cc3f0f0")
port map (
combout => N_52693,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03f3303ffc0ccfc0")
port map (
combout => N_53423,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03fc30cff30c3fc0")
port map (
combout => N_52716,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30cf03fc3fc0f30c")
port map (
combout => N_52739,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03fc30cff30c3fc0")
port map (
combout => N_52762,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30cf03fc3fc0f30c")
port map (
combout => N_52785,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0fc33c3cc3f0f0")
port map (
combout => N_52808,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0fc33c3cc3f0f0")
port map (
combout => N_52831,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_52854,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_52877,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_52900,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_52923,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_53441,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03fcf30c30cf3fc0")
port map (
combout => N_52946,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fccf00f33f0cc")
port map (
combout => N_52969,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fccf00f33f0cc")
port map (
combout => N_52992,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30cf3fc003fcf30c")
port map (
combout => N_52325,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_52348,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03fcf30c30cf3fc0")
port map (
combout => N_52371,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30cf3fc003fcf30c")
port map (
combout => N_52394,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_52417,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03fcf30c30cf3fc0")
port map (
combout => N_52440,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30cf3fc003fcf30c")
port map (
combout => N_52463,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_53464,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03fcf30c30cf3fc0")
port map (
combout => N_52486,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"303f03f3cfc0fc0c")
port map (
combout => N_52509,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c03f3fc3fcfc030")
port map (
combout => N_52532,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03fcf30c30cf3fc0")
port map (
combout => N_52555,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fccf00f33f0cc")
port map (
combout => N_52578,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33f0cc330fccf0")
port map (
combout => N_52601,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fccf00f33f0cc")
port map (
combout => N_52624,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fccf00f33f0cc")
port map (
combout => N_52647,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fccf00f33f0cc")
port map (
combout => N_52279,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fccf00f33f0cc")
port map (
combout => N_52302,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3003cffc3ff3c00c")
port map (
combout => N_53487,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33f0cc330fccf0")
port map (
combout => N_53510,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fccf00f33f0cc")
port map (
combout => N_53533,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fccf00f33f0cc")
port map (
combout => N_53015,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ffc33c3cc3ff00")
port map (
combout => N_53060,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0330fccff33f0cc0")
port map (
combout => N_53083,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_53106,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30033ff3cffcc00c")
port map (
combout => N_53129,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c33cffff3cc300")
port map (
combout => N_53152,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_6_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000c000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1685\,
dataf => N_32844_2,
datae => N_28681_I,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_27_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f003f00")
port map (
combout => N_33644,
dataf => N_33548,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_603\,
datad => N_33340_I,
datac => N_33178,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_12_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1633\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_O2_12_4\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(237));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_O2_25_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000ff000330ff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_875\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_I_O2_3_0\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff30000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_17\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_10\,
datae => N_28264_1,
datad => N_33735_1,
datac => N_34107,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0_O2_23_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff000c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8764\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8666\,
datae => N_32844_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11641\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
datab => N_34263_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_44_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_44__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8556\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_44__G2_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9486\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_1_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0330000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1187\,
dataf => N_33074_1,
datae => N_33652_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffa8aa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_16\,
dataf => N_33647,
datae => N_33655,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datac => N_33436_1,
datab => N_29071_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_34_0\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_31_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c300000000000000")
port map (
combout => N_33360,
dataf => N_28271_1,
datae => N_33144_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A21_1_RNI4GJF_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000f0c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
datad => N_32723_1,
datac => N_33340_I,
datab => N_28492_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_0_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000c300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9665\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
datad => N_34329_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9062\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8631\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9486\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_52288,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33330ff0ccccf0")
port map (
combout => N_52311,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03f3303ffc0ccfc0")
port map (
combout => N_52817,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"303f03f3cfc0fc0c")
port map (
combout => N_52518,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03f3303ffc0ccfc0")
port map (
combout => N_52771,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"303f03f3cfc0fc0c")
port map (
combout => N_53253,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"303f03f3cfc0fc0c")
port map (
combout => N_53184,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c3f03cff3c0fc30")
port map (
combout => N_52702,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c3f03cff3c0fc30")
port map (
combout => N_52886,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c3f03cff3c0fc30")
port map (
combout => N_52403,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"303f03f3cfc0fc0c")
port map (
combout => N_53092,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03f3303ffc0ccfc0")
port map (
combout => N_52610,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03f3303ffc0ccfc0")
port map (
combout => N_53001,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_53450,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03f3303ffc0ccfc0")
port map (
combout => N_53230,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03f3303ffc0ccfc0")
port map (
combout => N_53276,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"303f03f3cfc0fc0c")
port map (
combout => N_53299,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c3f03cff3c0fc30")
port map (
combout => N_53322,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c3f03cff3c0fc30")
port map (
combout => N_53345,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c3f03cff3c0fc30")
port map (
combout => N_52679,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c3f03cff3c0fc30")
port map (
combout => N_52725,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c3f03cff3c0fc30")
port map (
combout => N_52748,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33330ff0ccccf0")
port map (
combout => N_53473,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"303f03f3cfc0fc0c")
port map (
combout => N_52794,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"303f03f3cfc0fc0c")
port map (
combout => N_52840,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c3f03cff3c0fc30")
port map (
combout => N_52863,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c3f03cff3c0fc30")
port map (
combout => N_52909,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c3f03cff3c0fc30")
port map (
combout => N_52932,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c3f03cff3c0fc30")
port map (
combout => N_52955,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c3f03cff3c0fc30")
port map (
combout => N_52978,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_53496,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_52334,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_52357,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"303f03f3cfc0fc0c")
port map (
combout => N_52380,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03f3303ffc0ccfc0")
port map (
combout => N_52426,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"303f03f3cfc0fc0c")
port map (
combout => N_52449,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c3f03cff3c0fc30")
port map (
combout => N_52472,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03f3303ffc0ccfc0")
port map (
combout => N_52495,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_53069,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03f3303ffc0ccfc0")
port map (
combout => N_52541,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_52564,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"303f03f3cfc0fc0c")
port map (
combout => N_52587,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_52633,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33330ff0ccccf0")
port map (
combout => N_52656,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_53519,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_53542,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33330ff0ccccf0")
port map (
combout => N_53024,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_53049,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c3f03cff3c0fc30")
port map (
combout => N_53115,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03f3303ffc0ccfc0")
port map (
combout => N_53138,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_53161,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c3f03cff3c0fc30")
port map (
combout => N_53207,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_NOINSTANDNOEXC_0_A2_0_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cf00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_877_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1758\,
datae => N_33138_1,
datad => N_33607_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(66),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(67));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN18_LOCOV_RNIDLMG: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0fffffff3fff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_D\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5335\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(12),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.REEXCOVUV.UN13_LOCOV_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.REEXCOVUV.UN13_LOCOV_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_28_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1636\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_O2_10_4\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(250),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(254),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(255),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(256));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ffffccf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(19),
dataf => N_53931,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_21_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(21),
dataf => N_53930,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c0f00000c0c00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_4\,
dataf => N_32738_1,
datae => N_32844_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
datac => N_34341_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1749\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc00cc00f0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_1\,
dataf => N_32844_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9509\,
datad => N_34329_1,
datac => N_33607_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9566\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A26_12_0_RNIDE894_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffc0c0c0c0c0c0c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3945_I_I_O2_3_0\,
dataf => N_33070_1,
datae => N_34263_2,
datad => N_28857_1,
datac => N_28564_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A26_12_0\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1191\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datad => N_34263_2,
datac => N_28857_1,
datab => N_28266_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f3003300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1079\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11641\,
datae => N_33074_1,
datad => N_32782_1,
datac => N_34263_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_473\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O25_11_RNIRMPHE_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff000000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11641\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_782\,
datac => N_32782_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_604\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_3_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0003000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1048\,
dataf => N_32844_2,
datae => N_33070_1,
datad => N_33984_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_2_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000033303030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1647\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11641\,
datae => N_33340_I,
datad => N_28492_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9490\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1233\,
dataf => N_33074_1,
datae => N_33138_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_53016,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_53424,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff03c3c3c3c0ff0")
port map (
combout => N_53199,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30cf3fc003fcf30c")
port map (
combout => N_53222,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03fcf30c30cf3fc0")
port map (
combout => N_53245,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30cf3fc003fcf30c")
port map (
combout => N_53268,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_53291,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_53314,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_53337,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_52671,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_52694,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_52717,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff033cc33cc0ff0")
port map (
combout => N_53442,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03fcf30c30cf3fc0")
port map (
combout => N_52740,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30cf3fc003fcf30c")
port map (
combout => N_52763,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03fcf30c30cf3fc0")
port map (
combout => N_52786,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30cf3fc003fcf30c")
port map (
combout => N_52809,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_52832,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_52855,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_52878,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_52901,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_52924,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_52947,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_53465,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03fcf30c30cf3fc0")
port map (
combout => N_52970,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fccf00f33f0cc")
port map (
combout => N_52993,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fccf00f33f0cc")
port map (
combout => N_52326,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30cf3fc003fcf30c")
port map (
combout => N_52349,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_52372,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03fcf30c30cf3fc0")
port map (
combout => N_52395,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30cf3fc003fcf30c")
port map (
combout => N_52418,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fc33cf00f3cc3f0")
port map (
combout => N_52441,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03fcf30c30cf3fc0")
port map (
combout => N_52464,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30cf3fc003fcf30c")
port map (
combout => N_52487,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_53488,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03fcf30c30cf3fc0")
port map (
combout => N_52510,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c3c0ff00ff03c3c")
port map (
combout => N_52533,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c0f3cf00f3cf03c")
port map (
combout => N_52556,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3cf03c3c0f3cf0")
port map (
combout => N_52579,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_52602,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff033cc33cc0ff0")
port map (
combout => N_52625,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_52648,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_52280,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_52303,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_53511,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c0f3cf00f3cf03c")
port map (
combout => N_53061,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff033cc33cc0ff0")
port map (
combout => N_53534,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_53045,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33c33ccc333cc3cc")
port map (
combout => N_53084,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3cf03c3c0f3cf0")
port map (
combout => N_53107,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_53130,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c3c0ff00ff03c3c")
port map (
combout => N_53153,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c3c33cc33cc3c3c")
port map (
combout => N_53176,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_5_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc30cc0003cf33ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10875\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0c000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2_0\,
datae => N_32844_2,
datad => N_33070_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
datab => N_34341_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff5000dccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_10\,
dataf => N_33363,
datae => N_33548,
datad => N_33340_I,
datac => N_28564_2,
datab => N_33373_2,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_4_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000c000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9608\,
dataf => N_28264_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_43_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(43),
dataf => N_53880,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNINFNN_71_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcfffcfffcfff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(71));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_74_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0f0f0f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7274\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(62));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_M2_E: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0000000fc000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1028\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\,
datae => N_28857_1,
datad => N_33138_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9509\,
datab => N_32738_1_0);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_5_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0330000000000000")
port map (
combout => N_33027,
dataf => N_32909_1,
datae => N_29195_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(36),
dataf => N_53887,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff03ff0003030000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_584\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9486\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1586\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9502\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O17_3_RNIDGAND_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"44440000f444f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_7\,
dataf => N_33548,
datae => N_32723_1,
datad => N_33140_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_5_TZ\,
datab => N_33276,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A32_1_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000c0c0c000")
port map (
combout => N_33125,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_797\,
datae => N_32723_1,
datad => N_32796_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(18),
dataf => N_53923,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18));
\GRLFPC2_0_COMB_V_FSR_FCC_1_1_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc30ff00ff00ff00")
port map (
combout => \GRLFPC2_0.N_3226\,
dataf => \GRLFPC2_0.R.X.LD\,
datae => \GRLFPC2_0.R.X.AFSR\,
datad => CPO_CCZ(0),
datac => N_376,
datab => \GRLFPC2_0.N_1105\);
\GRLFPC2_0_COMB_V_FSR_FCC_1_1_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc30ff00ff00ff00")
port map (
combout => \GRLFPC2_0.N_3227\,
dataf => \GRLFPC2_0.R.X.LD\,
datae => \GRLFPC2_0.R.X.AFSR\,
datad => CPO_CCZ(1),
datac => N_377,
datab => \GRLFPC2_0.N_1105\);
GRLFPC2_0_V_FSR_AEXC_2_SQMUXA: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000c0f0f0f")
port map (
combout => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA\,
dataf => \GRLFPC2_0.N_1439\,
datae => \GRLFPC2_0.R.X.LD\,
datad => \GRLFPC2_0.R.X.AFSR\,
datac => \GRLFPC2_0.N_1517\,
datab => \GRLFPC2_0.N_1105\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_17_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => N_33913,
dataf => N_33735_1,
datae => N_32727_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_2_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1030\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datae => N_33340_I,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(42),
dataf => N_53919,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_7_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000030000000")
port map (
combout => N_33506,
dataf => N_28264_1,
datae => N_32796_2,
datad => N_28250_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_4_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000c0")
port map (
combout => N_34259,
dataf => N_33055,
datae => N_29071_1,
datad => N_33144_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000c00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1038\,
dataf => N_28857_1,
datae => N_28681_I,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0_O2_43_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000f000fcccf000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8556\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9525\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1586\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9514\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000300033003000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datae => N_34329_1,
datad => N_33507_1,
datac => N_33988_4,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff3000ba00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_9\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_603\,
datad => N_33574_1,
datac => N_28492_1,
datab => N_33179,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A32_2_0\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f333f000f000f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_3\,
dataf => N_33070_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9525\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9523\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1800\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffccf00000ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(34),
dataf => N_53889,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ffffccf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(38),
dataf => N_53919,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0002")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_6\,
dataf => N_34327,
datae => N_34333,
datad => N_33543,
datac => N_33721_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_604\,
dataa => N_34326_2);
GRLFPC2_0_R_I_RDD_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000fc30ff00")
port map (
combout => N_37429,
dataf => \GRLFPC2_0.N_1438_15\,
datae => \GRLFPC2_0.R.X.FPOP\,
datad => \GRLFPC2_0.R.I.RDD\,
datac => \GRLFPC2_0.R.X.RDD\,
datab => \GRLFPC2_0.N_1105\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f333f000f000f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_23\,
dataf => N_32738_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1595\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9598\,
datac => N_28390_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_3_S_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_A2_3_S\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1769\,
datad => N_32738_1_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datab => N_59);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_2_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"003c000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1082\,
dataf => N_33070_1,
datae => N_28312_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffccf00000ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(53),
dataf => N_53911,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_2_35_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000030000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9201\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datae => N_33074_1,
datad => N_34341_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_1_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c0000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1234\,
dataf => N_32782_1,
datae => N_34329_1,
datad => N_32722_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_4_1_RNIUTN28_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff73000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_0\,
datae => N_33070_1,
datad => N_33138_1,
datac => N_32859_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffcd000500")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_14\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_6\,
datae => N_32909_1,
datad => N_28212_1_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_604\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A32_13_1_0\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f888888888888888")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_0\,
dataf => N_33436_1,
datae => N_29195_1,
datad => N_32738_2,
datac => N_28549_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A11_3_1\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A11_3_0\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ffffccf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(55),
dataf => N_53914,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff04")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_20\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_14\,
datae => N_33225,
datad => N_33219,
datac => N_33548,
datab => N_28211_1,
dataa => N_33193);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_16_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"1300130013005f00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_16\(60),
dataf => N_28264_1,
datae => N_33074_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_0\(60),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_3_0\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A28_4_1\(60),
dataa => N_33710);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_24_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000c00000")
port map (
combout => N_34279,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11641\,
datae => N_32786_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00f000f3")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11641\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_571\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1607\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_30_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccfffff0cc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(30),
dataf => N_53889,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffeac0aa00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_9\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_4\,
datae => N_33138_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_13_0\(51),
datac => N_33577_1,
datab => N_34339_3,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_13_1\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ffffccf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(49),
dataf => N_53911,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff80")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_18\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_4\,
datae => N_34127,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_3\,
datac => N_32909_1,
datab => N_32786_1,
dataa => N_34256_1);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33c33ccc333cc3cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3c3c0ff03c3cf0")
port map (
combout => N_53146,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c0f0f3c3cf0f03c")
port map (
combout => N_53169,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3c3c0ff03c3cf0")
port map (
combout => N_53192,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c0f0f3c3cf0f03c")
port map (
combout => N_53215,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333c33c3cc3cccc")
port map (
combout => N_53238,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333c33c3cc3cccc")
port map (
combout => N_53261,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333c33c3cc3cccc")
port map (
combout => N_53284,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333c33c3cc3cccc")
port map (
combout => N_53307,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333c33c3cc3cccc")
port map (
combout => N_53330,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333c33c3cc3cccc")
port map (
combout => N_52664,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3cf03c3c0f3cf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3c3c0ff03c3cf0")
port map (
combout => N_52687,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c0f0f3c3cf0f03c")
port map (
combout => N_52710,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3c3c0ff03c3cf0")
port map (
combout => N_52733,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c0f0f3c3cf0f03c")
port map (
combout => N_52756,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333c33c3cc3cccc")
port map (
combout => N_52779,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333c33c3cc3cccc")
port map (
combout => N_52802,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333c33c3cc3cccc")
port map (
combout => N_52825,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33c33ccc333cc3cc")
port map (
combout => N_52848,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33c33ccc333cc3cc")
port map (
combout => N_52871,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33c33ccc333cc3cc")
port map (
combout => N_52894,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_53417,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3cf03c3c0f3cf0")
port map (
combout => N_52917,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_52940,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_52963,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c3c0ff00ff03c3c")
port map (
combout => N_52986,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c3c33cc33cc3c3c")
port map (
combout => N_52319,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff03c3c3c3c0ff0")
port map (
combout => N_52342,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c3c0ff00ff03c3c")
port map (
combout => N_52365,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c3c33cc33cc3c3c")
port map (
combout => N_52388,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff03c3c3c3c0ff0")
port map (
combout => N_52411,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c3c0ff00ff03c3c")
port map (
combout => N_52434,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_53435,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff03c3c3c3c0ff0")
port map (
combout => N_52457,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c3c0ff00ff03c3c")
port map (
combout => N_52480,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c333ccc333ccc3c")
port map (
combout => N_52503,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03f3303ffc0ccfc0")
port map (
combout => N_52526,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_52549,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33330ff0ccccf0")
port map (
combout => N_52572,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_52595,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_52618,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_52641,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_52273,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c0f0f3c3cf0f03c")
port map (
combout => N_53458,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33330ff0ccccf0")
port map (
combout => N_52296,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_53504,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_53527,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_53009,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330f0f33ccf0f0cc")
port map (
combout => N_53034,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333c33c3cc3cccc")
port map (
combout => N_53481,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3c3c0ff03c3cf0")
port map (
combout => N_53054,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33cc0ff00ff033cc")
port map (
combout => N_53077,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c0f0f3c3cf0f03c")
port map (
combout => N_53100,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333c33c3cc3cccc")
port map (
combout => N_53123,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00300000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_2\,
dataf => N_34194,
datae => N_32861_1,
datad => N_33340_I,
datac => N_33146_1,
datab => N_28564_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_10_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff000000ff404040")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_10\,
dataf => N_34029,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_4_1\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_4_0\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_6_1\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00fc000000f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_2\,
dataf => N_33070_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11641\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9522\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1713\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_17\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_10_0\,
datae => N_32899,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11641\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_525\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1044\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9486\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11641\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\,
datac => N_28857_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(47),
dataf => N_53901,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_9_I_O2_RNI678I3_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"303030fc000000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19\(9),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9486\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_525\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\,
datac => N_28266_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f333f000f000f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2_0\,
dataf => N_28266_2,
datae => N_28312_1,
datad => N_34133_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9511\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9368\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\,
datae => N_34329_1,
datad => N_29366_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0_O2_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000c0c0ccc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8631\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\,
datae => N_33340_I,
datad => N_28222_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9522\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_1_1_RNIFOC69_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff33000f00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_13_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_8\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\,
datad => N_34040_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_0_RNIDSOBU_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff00c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_17\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_13_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_9\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_13_TZ\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0800")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_8\,
dataf => N_32794,
datae => N_32792,
datad => N_29262_1,
datac => N_33297_1,
datab => N_33734_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff4000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_11\,
dataf => N_33911,
datae => N_33903,
datad => N_32738_1,
datac => N_33870,
datab => N_33734_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_17_RNIO51U3_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0200")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_3\,
datae => N_33588,
datad => N_28271_1,
datac => N_33178,
datab => N_28681_I,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"a0e4a0a000cc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_797\,
datae => N_28492_1,
datad => N_33111,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_9_0_0\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff3000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_21\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_17\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_9\,
datad => N_32908_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A32_0\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_0_RNIKHF73_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3f03300f0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_16__G2_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9522\,
datae => N_33369_1,
datad => N_32908_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0_0\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_15\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_8\,
datae => N_32738_1,
datad => N_29262_1,
datac => N_32723_1,
datab => N_28266_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff44004000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_3\,
dataf => N_33210,
datae => N_29653_1,
datad => N_28271_1,
datac => N_28227_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff1b000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_0\,
dataf => N_32916,
datae => N_32786_1,
datad => N_28251_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_9_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0f8f0088")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_8\,
dataf => N_34111,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_1_1\(54),
datad => N_34029,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_531\,
datab => N_33447_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_12_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aa00eac00000c0c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_603\,
datae => N_34329_1,
datad => N_33140_1,
datac => N_29366_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A32_11_0\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7_0\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_29_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000c000000000")
port map (
combout => N_33431,
dataf => N_33652_1,
datae => N_34341_1,
datad => N_33140_1,
datac => N_33146_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00000c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_13\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_719\,
datad => N_33146_1,
datac => N_28250_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff20")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_10_0\,
dataf => N_32908,
datae => N_32915,
datad => N_32917,
datac => N_34263_2,
datab => N_33436_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_33_0\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A28_2_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3000000f0000000")
port map (
combout => N_33721,
dataf => N_28266_2,
datae => N_33721_1,
datad => N_28261_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_0_A2_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000300000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_513\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_479\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f6f0f0f066000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A11_5_3\(61),
datae => N_33436_1,
datad => N_28208_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A11_5_2\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(33),
dataf => N_53896,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_17_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"135f5f5f00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_17\(60),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_11\(60),
datae => N_28264_1,
datad => N_33144_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A28_0_1\(60),
datab => N_33152_2,
dataa => N_33715);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff20")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_16_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_7\,
datae => N_33215,
datad => N_33220,
datac => N_32979_1,
datab => N_33178,
dataa => N_32722_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_0_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c300000000000000")
port map (
combout => N_32970,
dataf => N_34329_1,
datae => N_32722_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffccf00000ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(48),
dataf => N_53922,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ffffccf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(52),
dataf => N_53909,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_6_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => N_33028,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11641\,
datae => N_29262_1,
datad => N_33447_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O23_0_0_RNIMJ3M_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff00c8")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_10\,
dataf => N_33581,
datae => N_33574,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_782\,
datac => N_29071_1,
datab => N_32722_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_0_0\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ffffccf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(54),
dataf => N_53917,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_7_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf00c00030ff3ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10877\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff40")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_19\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_14\,
datae => N_34113,
datad => N_34114,
datac => N_33297_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_4_1\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f333f000f000f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_0\,
dataf => N_33507_1,
datae => N_33988_4,
datad => N_34047_2,
datac => N_34059_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffcf0eca0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_9\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9099\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9525\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1586\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9509\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1672\,
dataa => N_28390_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ff333cc0cc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(11),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(11),
datae => N_53929,
datad => N_53883,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_20_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(20),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(20),
datae => N_53923,
datad => N_53903,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_2_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0fcf0ff00cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9525\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1586\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9492\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9598\,
datab => N_32840_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff33300000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_769\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1647\,
datae => N_33070_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9525\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1800\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_O2_4_0_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000030ffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_O2_4_0\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1503\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_504\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1618\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_O2_12_RNI1QBR2_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fffcffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_4_TZ\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1852\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1503\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_504\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_9_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1519\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1497\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1496\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_451\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_504\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_I_A2_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000003000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1539\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1503\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_504\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1618\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_O2_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3f0330033003300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_544\,
dataf => N_32782_1,
datae => N_34341_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1595\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1592\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_812\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffc0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_1\,
dataf => N_34329,
datae => N_32818_I,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_3_0\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff8888888")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_7\,
dataf => N_34119,
datae => N_32909_1,
datad => N_33447_1,
datac => N_32818_I,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A24_0\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_15_0\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_1_A2_2_RNO_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fff0fcfffffffff")
port map (
combout => N_42365,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1633\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_446\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1637\,
datac => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(250));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_45_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1509\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1844\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_446\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(250));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_7_0_RNO_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fffffff0fcfffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_A2_7_8923_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_446\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1677\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1637\,
datac => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(250));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_2_RNII7LG_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff8")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_16\,
dataf => N_34059,
datae => N_34052,
datad => N_34041,
datac => N_34047,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9503\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9598\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff2")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9349\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_473\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9600\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_7_1_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"88cc88cc8888888c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_A2_7_1\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_473\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_661\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1809\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_479\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ff333cc0cc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(49),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(49),
datae => N_53888,
datad => N_53901,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_35_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff4")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_35__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8537\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9201\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9200\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9198\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9517\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_809\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_20_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cc00cc00fcf0cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_20__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_797\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9503\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9523\,
datac => N_33263_I,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1800\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_0_RNILQUF_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f30c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7035\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58));
\GRLFPC2_0_FPI_OP2_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(32),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_698,
datab => N_634);
\GRLFPC2_0_FPI_OP2_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(33),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_699,
datab => N_635);
\GRLFPC2_0_FPI_OP2_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(34),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_700,
datab => N_636);
\GRLFPC2_0_FPI_OP2_35_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(35),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_701,
datab => N_637);
\GRLFPC2_0_FPI_OP2_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(36),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_702,
datab => N_638);
\GRLFPC2_0_FPI_OP2_37_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(37),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_703,
datab => N_639);
\GRLFPC2_0_FPI_OP2_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(38),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_704,
datab => N_640);
\GRLFPC2_0_FPI_OP2_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(39),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_705,
datab => N_641);
\GRLFPC2_0_FPI_OP2_40_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(40),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_706,
datab => N_642);
\GRLFPC2_0_FPI_OP2_41_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(41),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_707,
datab => N_643);
\GRLFPC2_0_FPI_OP2_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(42),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_708,
datab => N_644);
\GRLFPC2_0_FPI_OP2_43_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(43),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_709,
datab => N_645);
\GRLFPC2_0_FPI_OP2_44_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(44),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_710,
datab => N_646);
\GRLFPC2_0_FPI_OP2_45_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(45),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_711,
datab => N_647);
\GRLFPC2_0_FPI_OP2_46_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(46),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_712,
datab => N_648);
\GRLFPC2_0_FPI_OP2_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(47),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_713,
datab => N_649);
\GRLFPC2_0_FPI_OP2_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(48),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_714,
datab => N_650);
\GRLFPC2_0_FPI_OP2_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(49),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_715,
datab => N_651);
\GRLFPC2_0_FPI_OP2_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(50),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_716,
datab => N_652);
\GRLFPC2_0_FPI_OP2_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(51),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_717,
datab => N_653);
\GRLFPC2_0_FPI_OP2_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(52),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_718,
datab => N_654);
\GRLFPC2_0_FPI_OP2_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(53),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_719,
datab => N_655);
\GRLFPC2_0_FPI_OP2_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(54),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_720,
datab => N_656);
\GRLFPC2_0_FPI_OP2_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(55),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_721,
datab => N_657);
\GRLFPC2_0_FPI_OP2_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(56),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_722,
datab => N_658);
\GRLFPC2_0_FPI_OP2_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(57),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_723,
datab => N_659);
\GRLFPC2_0_FPI_OP2_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(58),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_724,
datab => N_660);
\GRLFPC2_0_FPI_OP2_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(59),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_725,
datab => N_661);
\GRLFPC2_0_FPI_OP2_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(60),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_726,
datab => N_662);
\GRLFPC2_0_FPI_OP2_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(61),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_727,
datab => N_663);
\GRLFPC2_0_FPI_OP2_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(62),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_728,
datab => N_664);
\GRLFPC2_0_FPI_OP2_63_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP2\(63),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\,
datac => N_729,
datab => N_665);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_3_RNI771D2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c0ff3fff3f00c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_116\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_60.Z_1_CO1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_3_RNI771D2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00c000c00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_319__G1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_116\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_60.Z_1_CO1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7045\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7038\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2_3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_13\,
dataf => N_33646,
datae => N_33648,
datad => N_32861_1,
datac => N_32982_1,
datab => N_29366_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(38),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(38),
datae => N_53887,
datad => N_53885,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_20_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0015000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_20\(60),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_5\(60),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_6\(60),
datad => N_33721,
datac => N_28264_1,
datab => N_33735_3,
dataa => N_34268);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_22\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_7\,
datad => N_33650,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_8_1\,
datab => N_33643,
dataa => N_33654);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffa0ec")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_20\,
dataf => N_33125,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_8\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
datac => N_33175,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A32_19_0\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_18_TZ\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_45_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9159\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8573\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2_1\,
datac => N_32762_I,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1736\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9479\);
\GRLFPC2_0_FPI_OP1_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP1\(32),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS1\(0),
datad => \GRLFPC2_0.R.A.RS1D\,
datac => N_666,
datab => N_602);
\GRLFPC2_0_FPI_OP1_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP1\(33),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS1\(0),
datad => \GRLFPC2_0.R.A.RS1D\,
datac => N_667,
datab => N_603);
\GRLFPC2_0_FPI_OP1_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP1\(34),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS1\(0),
datad => \GRLFPC2_0.R.A.RS1D\,
datac => N_668,
datab => N_604);
\GRLFPC2_0_FPI_OP1_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP1\(36),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS1\(0),
datad => \GRLFPC2_0.R.A.RS1D\,
datac => N_670,
datab => N_606);
\GRLFPC2_0_FPI_OP1_37_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP1\(37),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS1\(0),
datad => \GRLFPC2_0.R.A.RS1D\,
datac => N_671,
datab => N_607);
\GRLFPC2_0_FPI_OP1_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP1\(38),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS1\(0),
datad => \GRLFPC2_0.R.A.RS1D\,
datac => N_672,
datab => N_608);
\GRLFPC2_0_FPI_OP1_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP1\(39),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS1\(0),
datad => \GRLFPC2_0.R.A.RS1D\,
datac => N_673,
datab => N_609);
\GRLFPC2_0_FPI_OP1_41_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP1\(41),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS1\(0),
datad => \GRLFPC2_0.R.A.RS1D\,
datac => N_675,
datab => N_611);
\GRLFPC2_0_FPI_OP1_43_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP1\(43),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS1\(0),
datad => \GRLFPC2_0.R.A.RS1D\,
datac => N_677,
datab => N_613);
\GRLFPC2_0_FPI_OP1_44_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP1\(44),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS1\(0),
datad => \GRLFPC2_0.R.A.RS1D\,
datac => N_678,
datab => N_614);
\GRLFPC2_0_FPI_OP1_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP1\(47),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS1\(0),
datad => \GRLFPC2_0.R.A.RS1D\,
datac => N_681,
datab => N_617);
\GRLFPC2_0_FPI_OP1_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP1\(49),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS1\(0),
datad => \GRLFPC2_0.R.A.RS1D\,
datac => N_683,
datab => N_619);
\GRLFPC2_0_FPI_OP1_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP1\(51),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS1\(0),
datad => \GRLFPC2_0.R.A.RS1D\,
datac => N_685,
datab => N_621);
\GRLFPC2_0_FPI_OP1_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP1\(53),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS1\(0),
datad => \GRLFPC2_0.R.A.RS1D\,
datac => N_687,
datab => N_623);
\GRLFPC2_0_FPI_OP1_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP1\(54),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS1\(0),
datad => \GRLFPC2_0.R.A.RS1D\,
datac => N_688,
datab => N_624);
\GRLFPC2_0_FPI_OP1_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP1\(55),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS1\(0),
datad => \GRLFPC2_0.R.A.RS1D\,
datac => N_689,
datab => N_625);
\GRLFPC2_0_FPI_OP1_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP1\(56),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS1\(0),
datad => \GRLFPC2_0.R.A.RS1D\,
datac => N_690,
datab => N_626);
\GRLFPC2_0_FPI_OP1_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP1\(57),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS1\(0),
datad => \GRLFPC2_0.R.A.RS1D\,
datac => N_691,
datab => N_627);
\GRLFPC2_0_FPI_OP1_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP1\(58),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS1\(0),
datad => \GRLFPC2_0.R.A.RS1D\,
datac => N_692,
datab => N_628);
\GRLFPC2_0_FPI_OP1_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP1\(59),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS1\(0),
datad => \GRLFPC2_0.R.A.RS1D\,
datac => N_693,
datab => N_629);
\GRLFPC2_0_FPI_OP1_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP1\(60),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS1\(0),
datad => \GRLFPC2_0.R.A.RS1D\,
datac => N_694,
datab => N_630);
\GRLFPC2_0_FPI_OP1_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP1\(61),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS1\(0),
datad => \GRLFPC2_0.R.A.RS1D\,
datac => N_695,
datab => N_631);
\GRLFPC2_0_FPI_OP1_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.FPI.OP1\(62),
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS1\(0),
datad => \GRLFPC2_0.R.A.RS1D\,
datac => N_696,
datab => N_632);
\GRLFPC2_0_FPI_OP1_I_M3_45_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0ccf0cccc")
port map (
combout => \GRLFPC2_0.N_71\,
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS1\(0),
datad => \GRLFPC2_0.R.A.RS1D\,
datac => N_679,
datab => N_615);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c0c0c0c0eaeaeac0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_11_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_797\,
datae => N_33543,
datad => N_28212_1_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_11_0\(51),
datab => N_33738_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A21_0\(51));
\GRLFPC2_0_R_A_RF2REN_RNO_0_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00fc000000ff00ff")
port map (
combout => N_37387,
dataf => \GRLFPC2_0.N_1714_I\,
datae => \GRLFPC2_0.N_1093\,
datad => \GRLFPC2_0.N_1072\,
datac => \GRLFPC2_0.COMB.FPDECODE.ST\,
datab => \GRLFPC2_0.N_951\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_30_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffdc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_30__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_759\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_769\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_30__G2_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1832\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_30__G2_1\,
dataa => N_28261_1);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_3_RNIM0F91_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00c000c00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_959_I\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_57\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_1_CO0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_3_RNIM0F91: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c0ff3fff3f00c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SBLSBS_2\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_57\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_1_CO0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_0_37_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff8888888")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_756\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1718\,
datae => N_32738_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9486\,
datac => N_32782_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9502\,
dataa => N_28390_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_0_0_RNID0KJ3_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffa7700f7f07700")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_11\,
dataf => N_32727_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_0_0\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_2_0\(31),
datac => N_33985_2,
datab => N_33560,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffc0c0c0c0c0c0c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_1\,
dataf => N_32738_1,
datae => N_28266_2,
datad => N_32840_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9514\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9570\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_0_RNI3O5P_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff1000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9371\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9369\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9486\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8619\,
dataa => N_34326_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_3_RNISQCT_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1048\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9375\,
datac => N_33735_1,
datab => N_33146_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9490\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_13\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_1\,
datae => N_33830,
datad => N_33842,
datac => N_33832,
datab => N_33844,
dataa => N_33845);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_13_RNIS7OJ3_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffff8f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_12\,
dataf => N_33572,
datae => N_33576,
datad => N_32730_1,
datac => N_33584,
datab => N_33565,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(55),
datae => N_53911,
datad => N_53913,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000f888")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_9\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1200\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datad => N_28857_1,
datac => N_28266_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1595\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_0_RNI7LUH3_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff0c00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_6\,
dataf => N_34039,
datae => N_33447_1,
datad => N_28261_1,
datac => N_34132_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_35_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(35),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(35),
datae => N_53896,
datad => N_53904,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff8888888f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_473\,
datad => N_34029,
datac => N_33146_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1595\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9547\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_39__G2_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1135\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1134\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1133\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_525\,
datab => N_32782_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_37_1_RNIRG6F8_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffce")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_18\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_8\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_10\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_11\,
datac => N_33548,
datab => N_33590,
dataa => N_33373_2);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_MIFROMINST: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c400c4c4cc00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3924\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1758\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_473\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.MIFROMINST_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(63));
GRLFPC2_0_COMB_V_I_RDD_1_I_A3_15_RNIHJLA: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffff000000")
port map (
combout => \GRLFPC2_0.N_1876_2\,
dataf => \GRLFPC2_0.N_54\,
datae => \GRLFPC2_0.N_1438_15\,
datad => N_13);
\GRLFPC2_0_R_I_EXC_RNO_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00030000000f0000")
port map (
combout => \GRLFPC2_0.R.I.EXC_2_0_3__G2\,
dataf => \GRLFPC2_0.N_1438_15\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(40),
datab => N_13);
GRLFPC2_0_R_I_V_ENA_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00cc000c")
port map (
combout => \GRLFPC2_0.R.I.V_1_0_G2\,
dataf => \GRLFPC2_0.N_54\,
datae => \GRLFPC2_0.N_1438_15\,
datad => \GRLFPC2_0.COMB.ANNULRES_1\,
datac => N_13,
datab => N_11);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_759\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1648\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9600\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_493\);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_23_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0ff00cccc")
port map (
combout => \GRLFPC2_0.N_3106\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.FSR.TEM\(0),
datac => N_689,
datab => N_625);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcf3f00f0c0300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(38),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(37),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ff0f0f3333")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(49),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_71_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00030000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.UN36_PCTRL_NEW_I\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3924\,
datae => \GRLFPC2_0.N_3475\,
datad => \GRLFPC2_0.R.MK.RST\,
datac => \GRLFPC2_0.N_67\,
datab => \GRLFPC2_0.R.MK.RST2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccfff0ffcc00f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(29),
dataf => N_53969,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_6_1_RNI057G3_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffd5c0c0c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_7\,
dataf => N_33589,
datae => N_33652_1,
datad => N_29071_1,
datac => N_29366_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_6_1\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_45_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ffcc00f000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(45),
dataf => N_53973,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0ff00cccc")
port map (
combout => \GRLFPC2_0.N_3090\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.FSR.AEXC\(2),
datac => N_673,
datab => N_609);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_82_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0ff00ccccff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(82),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => N_696,
datac => N_667,
datab => N_603);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf3f0ff0c03000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(56),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(56),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0ff00ccccff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(83),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => N_695,
datac => N_666,
datab => N_602);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff33ffffff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ffcc00f000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(38),
dataf => N_53988,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_16_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ffcc00f000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(16),
dataf => \GRLFPC2_0.FPI.OP2\(41),
datae => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_704,
datab => N_640);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0ff00cccc")
port map (
combout => \GRLFPC2_0.N_3108\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.FSR.TEM\(2),
datac => N_691,
datab => N_627);
\GRLFPC2_0_R_FSR_FTT_RNO_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f0c000f000")
port map (
combout => \GRLFPC2_0.R.FSR.FTT_0_0_0__G1\,
dataf => \GRLFPC2_0.N_1015\,
datae => \GRLFPC2_0.N_58\,
datad => \GRLFPC2_0.R.FSR.FTT\(0),
datac => N_11,
datab => \GRLFPC2_0.N_1105\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000fc0000000c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10079\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9783\,
datae => \GRLFPC2_0.FPI.LDOP_1\,
datad => \GRLFPC2_0.FPI.RST_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(171));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000fc0000000c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10078\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9782\,
datae => \GRLFPC2_0.FPI.LDOP_1\,
datad => \GRLFPC2_0.FPI.RST_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(172));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000fc0000000c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10077\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9781\,
datae => \GRLFPC2_0.FPI.LDOP_1\,
datad => \GRLFPC2_0.FPI.RST_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(173));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0fcfffff0ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856\,
datae => \GRLFPC2_0.FPI.LDOP_1_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895\,
datac => \GRLFPC2_0.FPI.RST_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_RNIHQ2Q4_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300030303000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(58),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(58),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_317__G1\,
datac => \GRLFPC2_0.FPI.LDOP_1_2\,
datab => \GRLFPC2_0.FPI.RST_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9988\,
dataf => \GRLFPC2_0.FPI.LDOP_1_2\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(142),
datab => N_726);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9987\,
dataf => \GRLFPC2_0.FPI.LDOP_1_2\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(143),
datab => N_725);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9986\,
dataf => \GRLFPC2_0.FPI.LDOP_1_2\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(144),
datab => N_724);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9985\,
dataf => \GRLFPC2_0.FPI.LDOP_1_2\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(145),
datab => N_723);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_30_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9984\,
dataf => \GRLFPC2_0.FPI.LDOP_1_2\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(146),
datab => N_722);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9983\,
dataf => \GRLFPC2_0.FPI.LDOP_1_2\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(147),
datab => N_721);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9982\,
dataf => \GRLFPC2_0.FPI.LDOP_1_2\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(148),
datab => N_720);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9980\,
dataf => \GRLFPC2_0.FPI.LDOP_1_2\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(150),
datab => N_718);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_35_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9979\,
dataf => \GRLFPC2_0.FPI.LDOP_1_2\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(151),
datab => N_717);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9978\,
dataf => \GRLFPC2_0.FPI.LDOP_1_2\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(152),
datab => N_716);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_37_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9977\,
dataf => \GRLFPC2_0.FPI.LDOP_1_2\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(153),
datab => N_715);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9976\,
dataf => \GRLFPC2_0.FPI.LDOP_1_2\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(154),
datab => N_714);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9975\,
dataf => \GRLFPC2_0.FPI.LDOP_1_2\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(155),
datab => N_713);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_40_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9974\,
dataf => \GRLFPC2_0.FPI.LDOP_1_2\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(156),
datab => N_712);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_41_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9973\,
dataf => \GRLFPC2_0.FPI.LDOP_1\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(157),
datab => N_711);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9972\,
dataf => \GRLFPC2_0.FPI.LDOP_1\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(158),
datab => N_710);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_43_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9971\,
dataf => \GRLFPC2_0.FPI.LDOP_1\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(159),
datab => N_709);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_44_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9970\,
dataf => \GRLFPC2_0.FPI.LDOP_1\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(160),
datab => N_708);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_45_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9969\,
dataf => \GRLFPC2_0.FPI.LDOP_1\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(161),
datab => N_707);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_46_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9968\,
dataf => \GRLFPC2_0.FPI.LDOP_1\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(162),
datab => N_706);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9967\,
dataf => \GRLFPC2_0.FPI.LDOP_1\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(163),
datab => N_705);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9966\,
dataf => \GRLFPC2_0.FPI.LDOP_1\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(164),
datab => N_704);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9964\,
dataf => \GRLFPC2_0.FPI.LDOP_1\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(166),
datab => N_702);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9963\,
dataf => \GRLFPC2_0.FPI.LDOP_1\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(167),
datab => N_701);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9962\,
dataf => \GRLFPC2_0.FPI.LDOP_1\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(168),
datab => N_700);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9961\,
dataf => \GRLFPC2_0.FPI.LDOP_1\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(169),
datab => N_699);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc00cc00ccf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9960\,
dataf => \GRLFPC2_0.FPI.LDOP_1\,
datae => \GRLFPC2_0.FPI.RST_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(170),
datab => N_698);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_43_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ffcc00f000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(43),
dataf => N_53972,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_15_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ffcc00f000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(15),
dataf => N_53956,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1036\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1030\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1027\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_46_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ff0f0f3333")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(46),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0ff00cccc")
port map (
combout => \GRLFPC2_0.N_3109\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.FSR.TEM\(3),
datac => N_692,
datab => N_628);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_74_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0fff000ccffcc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(74),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.FPI.OP1\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_675,
datab => N_611);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0f0f00ff3333")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(48),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00ff0f0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(50),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_44_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ffccfff000cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(44),
dataf => N_53952,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ffccfff000cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(10),
dataf => N_53984,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_14_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ffcc00f000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(14),
dataf => N_53959,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff02")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1697\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1028\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_797\,
datab => N_33436_1,
dataa => N_32840_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ffccfff000cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(33),
dataf => N_53976,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_21_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccfff0ffcc00f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(21),
dataf => N_53979,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffccfff000cc00f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(25),
dataf => N_53969,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0fff000ccffcc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(61),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.FPI.OP1\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_688,
datab => N_624);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffeac0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_11\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_8\,
datae => N_33661,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_52_0\(58),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_28_1\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_28_0\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_52_1\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_71_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0fff000ccffcc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(71),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.FPI.OP1\(41),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_678,
datab => N_614);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_78_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff000f0ffcc00cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(78),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.FPI.OP1\(37),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_668,
datab => N_604);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_81_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0ff00ccccff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(81),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => N_697,
datac => N_668,
datab => N_604);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_40_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ffcc00f000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(40),
dataf => N_53952,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff33ffffff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00ff0f0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(51),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_30_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ffccfff000cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(30),
dataf => N_53989,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ffcc00f000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(18),
dataf => \GRLFPC2_0.FPI.OP2\(39),
datae => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_702,
datab => N_638);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccfff0ffcc00f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(19),
dataf => N_53956,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_76_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff000f0ffcc00cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(76),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.FPI.OP1\(39),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_670,
datab => N_606);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_79_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0fff000ccffcc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(79),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.FPI.OP1\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_670,
datab => N_606);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3fcf00f030c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(52),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(51),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3fcf0ff030c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(53),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff3")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10195\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_21_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff000f0ffcc00cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(21),
dataf => \GRLFPC2_0.COMB.UN1_FPCI_4\,
datae => \GRLFPC2_0.FPI.OP2\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_699,
datab => N_635);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcf3f00f0c0300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(53),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf3f0ff0c03000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(55),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_68_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0fff000ccffcc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(68),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.FPI.OP1\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_681,
datab => N_617);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_240_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bb00ff00b800fc00")
port map (
combout => N_37419,
dataf => \GRLFPC2_0.FPO.EXP\(4),
datae => N_37019_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_240__G2_0_7674_I_0\,
datac => \GRLFPC2_0.FPI.LDOP_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(253));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_3_RNITBMG1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bb00ff00b800fc00")
port map (
combout => N_37418,
dataf => \GRLFPC2_0.FPO.EXP\(3),
datae => N_37019_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_241__G2_0_7643_I_0\,
datac => \GRLFPC2_0.FPI.LDOP_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(254));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CARRY_0_RNI15IF1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bb00ff00b800fc00")
port map (
combout => N_37415,
dataf => \GRLFPC2_0.FPO.EXP\(0),
datae => N_37019_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__G2_0_7550_I_0\,
datac => \GRLFPC2_0.FPI.LDOP_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(257));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_242_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bb00ff00b800fc00")
port map (
combout => N_37417,
dataf => \GRLFPC2_0.FPO.EXP\(2),
datae => N_37019_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_242__G2_0_7612_I_0\,
datac => \GRLFPC2_0.FPI.LDOP_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(255));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcff3c33c0c3000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(29),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(28),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"303000aafcfc00aa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10133\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
datad => \GRLFPC2_0.FPI.LDOP_0_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(117));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_248_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffaa303055003030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(248),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10512\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10530\,
datad => \GRLFPC2_0.FPO.EXP\(9),
datac => \GRLFPC2_0.FPI.OP1\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_16_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00fcfcff000c0c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10118\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9822\,
datae => \GRLFPC2_0.FPI.LDOP_0_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(132));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00fcfcff000c0c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10116\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9820\,
datae => \GRLFPC2_0.FPI.LDOP_0_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(134));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_21_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00fcfcff000c0c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10113\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9817\,
datae => \GRLFPC2_0.FPI.LDOP_0_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(137));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9166\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1212\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1214\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_797\,
datab => N_28681_I,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1714\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_CIN_1_RNI36L31: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccc3c333333c3ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_116\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58\(56),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1274_I\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_23_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff8")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_23__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8764\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1301\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1303\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1302\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9503\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9498\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_I_O2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffa000ffffeccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1846\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1539\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1852\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1839\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1618\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0800")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_14\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1191\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_12\,
datad => N_28634_1,
datac => N_33548,
datab => N_28658_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ffaafcfcffaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10132\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
datad => \GRLFPC2_0.FPI.LDOP_0_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(118));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_238_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bb00ff00b800fc00")
port map (
combout => N_37421,
dataf => \GRLFPC2_0.FPO.EXP\(6),
datae => N_37019_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_238__G2_0_7736_I_0\,
datac => \GRLFPC2_0.FPI.LDOP_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(251));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIRBMG1_256_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bb00ff00b800fc00")
port map (
combout => N_37416,
dataf => \GRLFPC2_0.FPO.EXP\(1),
datae => N_37019_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_243__G2_0_7581_I_0\,
datac => \GRLFPC2_0.FPI.LDOP_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(256));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0c00aafcfc00aa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10134\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
datad => \GRLFPC2_0.FPI.LDOP_0_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(116));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_10_RNI8SHT3_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff2")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_14\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9373\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1055\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_525\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9600\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_1_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffc0c0ffc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1082\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_525\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9600\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1592\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_4_0\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_8\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_758\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_7\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8573\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_237_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bb00ff00b800fc00")
port map (
combout => N_37422,
dataf => \GRLFPC2_0.FPO.EXP\(7),
datae => N_37019_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_237__G2_0_7767_I_0\,
datac => \GRLFPC2_0.FPI.LDOP_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(250));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_20\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_16\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_10\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_11\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_76_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333f333f333fffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7272\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_663\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_239_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"bb00ff00b800fc00")
port map (
combout => N_37420,
dataf => \GRLFPC2_0.FPO.EXP\(5),
datae => N_37019_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_239__G2_0_7705_I_0\,
datac => \GRLFPC2_0.FPI.LDOP_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(252));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"50fa51fb54fe55ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(6),
datad => N_54021,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_13\,
dataf => N_33916,
datae => N_33904,
datad => N_33895,
datac => N_33897);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_O2_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3f3f3f3f3333333")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_513\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_458\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_426\,
datad => N_32738_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(67),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(66));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_PCTRL_NEW_1_S: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000300000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_513\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_877_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_551\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_TEMP: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00c0ffff00cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856\,
datae => \GRLFPC2_0.FPI.LDOP_0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(21));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTABORTNULLEXC_RNIBVBO5: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cccc00c0cccc00cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856\,
datae => \GRLFPC2_0.FPI.LDOP_0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNI9VBO5_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cccc00c0cccc00cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856\,
datae => \GRLFPC2_0.FPI.LDOP_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3fcf0ff030c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(27),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(27),
datae => N_53969,
datad => N_53976,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00cfcfff000303")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(48),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(50),
datac => N_53953,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_PCTRL_1_CO3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_43_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3ffc0fff300c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(43),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(43),
datae => N_53971,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datac => N_53973,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"50fa51fb54fe55ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(32),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(31),
datad => N_54012,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN2_MIXOIN_1_RNI37AL7_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff9fef7f9fff7fe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SBLSBS_1\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SBLSBS_2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_959_I\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1_1\,
datab => N_53998,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5452\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000003000030033")
port map (
combout => N_54031,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_23_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcfffc0030ff3000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(23),
dataf => N_53969,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(23),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datac => N_53958,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIIGMJP_66_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff0f00000f0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_51_I\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_475\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(67),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(66));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_I_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00f0fffff0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_475\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(67),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(66));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffcff0f0f0c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10197\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(55),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf3f0ff0c03000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(38),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(38),
datae => N_53952,
datad => N_53961,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_U: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000d050f05")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR\,
dataf => N_53985,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23_1_SUM_0_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cc333cc33cc333cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1281_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7035\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7034\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_50_1_SUM_0_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cc333cc33cc333cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1281_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7035\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7051\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_1_A2_2_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cc00c00000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_A2_1_A2_2\(83),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_513\,
datae => N_28511,
datad => N_42365,
datac => N_28510,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1618\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNI5KFP5_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcfc0000fcfc00fc")
port map (
combout => N_61580,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_49_I\,
datae => \GRLFPC2_0.FPI.LDOP_0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_RNIPSLS5: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f3f0f3f0f3")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_49_I\,
datac => \GRLFPC2_0.FPI.LDOP_0_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNI9KFP5_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcfc0000fcfc0030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_49_I\,
datae => \GRLFPC2_0.FPI.LDOP_0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"5072d8fa5577ddff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(29),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(29),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(30),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_22_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"50d872fa55dd77ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(22),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(22),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(22),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNITKPG_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000fc00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10530\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\,
datad => \GRLFPC2_0.FPI.LDOP_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00fffcff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\,
datad => \GRLFPC2_0.FPI.LDOP_0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPBREGLOADEN: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00fffcff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\,
datad => \GRLFPC2_0.FPI.LDOP_0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_17_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f01000f0f0f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1540\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_386\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_893\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1636\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1618\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_I_O2_3_0\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"5072d8fa5577ddff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(26),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(26),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"5055d8dd7277faff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8_I\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_247_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30ff303030003030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(247),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10527\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
datad => \GRLFPC2_0.FPI.LDOP_0_0\,
datac => \GRLFPC2_0.FPI.OP1\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_249_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30ff303030003030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(249),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10525\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
datad => \GRLFPC2_0.FPI.LDOP_0_0\,
datac => \GRLFPC2_0.FPI.OP1\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_246_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fafa00cc505000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(246),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10514\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10530\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SS0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffff003f00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0_N_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0_M3_I_A3_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_9_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000effeffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_9\(47),
dataf => N_34257,
datae => N_34256_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_29_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3020000000000000")
port map (
combout => N_32907,
dataf => N_34263_2,
datae => N_33436_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_RESULT_IV_0_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"155515551555d555")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_0\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SFTLFT.AREGXORBREG\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_1_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0024000000000000")
port map (
combout => N_33500,
dataf => N_28271_1,
datae => N_33899_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_4_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c050000000000000")
port map (
combout => N_33288,
dataf => N_33138_1,
datae => N_32796_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_1_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"8ca0000000000000")
port map (
combout => N_33023,
dataf => N_29071_1,
datae => N_28492_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A24_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff3000000000000")
port map (
combout => N_34180,
dataf => N_28634_1,
datae => N_32731_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A15_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000232c0000")
port map (
combout => N_33021,
dataf => N_33004,
datae => N_33146_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_0_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cff0000000000000")
port map (
combout => N_33208,
dataf => N_32844_3,
datae => N_33503_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83));
GRLFPC2_0_COMB_V_A_SEQERR_1_0_O2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"2022c00c20222022")
port map (
combout => \GRLFPC2_0.N_94\,
dataf => \GRLFPC2_0.FPCI_O\(59),
datae => \GRLFPC2_0.FPCI_O\(58),
datad => \GRLFPC2_0.R.STATE_O\(0),
datac => \GRLFPC2_0.R.STATE_O\(1),
datab => \GRLFPC2_0.FPCI_O\(60),
dataa => \GRLFPC2_0.N_1837_O\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_0_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00220000a0a00000")
port map (
combout => N_33777,
dataf => N_33146_1,
datae => N_32738_2,
datad => N_28681_I,
datac => N_34254_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_13_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"033307770fff0fff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_13\(11),
dataf => N_33725_1,
datae => N_33507_1,
datad => N_28564_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A26_12_0\(11),
datab => N_28250_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf0cc00f0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_7\,
dataf => N_28634_1,
datae => N_28222_1,
datad => N_32727_1,
datac => N_33735_3,
datab => N_34055_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc50dc00cc00cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_1\,
dataf => N_33070_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_797\,
datac => N_33138_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1659\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_11_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000001000000000")
port map (
combout => N_33510,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_719\,
datae => N_33368_1,
datad => N_28211_1,
datac => N_32908_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_604\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_10_2_RNIFRK56_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccfccccc00f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_4\,
dataf => N_33794,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11641\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9503\,
datab => N_32732_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A8_4_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000200")
port map (
combout => N_28254,
dataf => N_32844_2,
datae => N_29653_1,
datad => N_34263_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_797\,
datab => N_28652_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A22_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ed00a50000000000")
port map (
combout => N_33827,
dataf => N_28560_2,
datae => N_33798_I,
datad => N_33734_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN11_WQSTSETS: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f7f7f707")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN11_WQSTSETS\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TEMP\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(14));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffc0c0c0c0c0c0c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_3\,
dataf => N_32738_1,
datae => N_29262_1,
datad => N_33447_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_15_1\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_15_0\(54));
GRLFPC2_0_R_FSR_NONSTD_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"b888b888fccc3000")
port map (
combout => \GRLFPC2_0.R.FSR.NONSTD_0_0_G1\,
dataf => \GRLFPC2_0.N_1171\,
datae => \GRLFPC2_0.R.FSR.NONSTD\,
datad => N_428,
datac => N_11,
datab => \GRLFPC2_0.N_3027\,
dataa => N_388);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_3_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0330000000000000")
port map (
combout => N_34114,
dataf => N_28264_1,
datae => N_32858_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_6_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0bbb0fffbbbbffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_6\(60),
dataf => N_33074_1,
datae => N_32982_1,
datad => N_28560_2,
datac => N_33756,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_13_1\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_12_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333ffffff3fffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_12\(11),
dataf => N_28634_1,
datae => N_34007,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_7_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000008800000")
port map (
combout => N_34118,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_603\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_531\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_6_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"007f7f7f00ffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_6\(11),
dataf => N_32861_1,
datae => N_33574_1,
datad => N_33985_2,
datac => N_33984_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_2_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"5450000000000000")
port map (
combout => N_33024,
dataf => N_33659_1,
datae => N_34329_1,
datad => N_29366_1,
datac => N_32738_1_0,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_8_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3033300000000000")
port map (
combout => N_34047,
dataf => N_34047_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83));
GRLFPC2_0_COMB_UN6_IUEXEC_I: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000200")
port map (
combout => \GRLFPC2_0.N_54\,
dataf => \GRLFPC2_0.R.MK.RST\,
datae => \GRLFPC2_0.N_1714_I\,
datad => \GRLFPC2_0.N_3545\,
datac => \GRLFPC2_0.R.MK.RST2\,
datab => \GRLFPC2_0.COMB.ANNULFPU_1_O_0\,
dataa => \GRLFPC2_0.R.MK.BUSY_O\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_6_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000030000000000")
port map (
combout => N_33505,
dataf => N_28271_1,
datae => N_33984_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_X2_RNIR9RQ_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"55d500c000c000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_3\,
dataf => N_28264_1,
datae => N_33070_1,
datad => N_33548,
datac => N_33503_1,
datab => N_28892_I,
dataa => N_33547_I);
\GRLFPC2_0_R_FSR_RD_RNO_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"b888b888fccc3000")
port map (
combout => \GRLFPC2_0.R.FSR.RD_0_0_0__G1\,
dataf => \GRLFPC2_0.N_1171\,
datae => \GRLFPC2_0.R.FSR.RD\(0),
datad => N_436,
datac => N_11,
datab => \GRLFPC2_0.N_3027\,
dataa => N_396);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_2_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"55ff45cfffffcfcf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_2\(47),
dataf => N_28264_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_782\,
datad => N_29071_1,
datac => N_32909_1,
datab => N_29195_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f7f7f0f0f777f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_10_TZ\,
dataf => N_33659_1,
datae => N_28634_1,
datad => N_28857_1,
datac => N_33144_1,
datab => N_33179,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_3_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"135fffff33ffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_3\(11),
dataf => N_33340_I,
datae => N_32786_1,
datad => N_28250_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A24_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c4c0000000000000")
port map (
combout => N_32777,
dataf => N_32861_1,
datae => N_32844_3,
datad => N_33984_2,
datac => N_33734_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"6eeaf7bffb7f9dd5")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5301\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5339\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10880\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10882\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A25_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ea000000000000")
port map (
combout => N_33351,
dataf => N_33074_1,
datae => N_28564_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_3_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3f773fffff77ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_3\(60),
dataf => N_29653_1,
datae => N_33735_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_531\,
datac => N_33081_1,
datab => N_28250_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_0_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30000000f000f000")
port map (
combout => N_33896,
dataf => N_33004,
datae => N_29195_1,
datad => N_33503_1,
datac => N_28921_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"8888a0000000a000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_3\,
dataf => N_32861_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_531\,
datad => N_33721_1,
datac => N_32859_1,
datab => N_28652_1,
dataa => N_28251_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A24_RNI7H967_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00009000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_0\,
dataf => N_34180,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\,
datad => N_28857_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcf00000cc000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_4\,
dataf => N_32861_1,
datae => N_28658_1,
datad => N_34335_2,
datac => N_34340_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"8004000000040000")
port map (
combout => N_34254,
dataf => N_32738_1,
datae => N_34254_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_5_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000088000000000")
port map (
combout => N_34330,
dataf => N_33652_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_531\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
\GRLFPC2_0_R_FSR_RD_RNO_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"b888b888fccc3000")
port map (
combout => \GRLFPC2_0.R.FSR.RD_0_0_1__G1\,
dataf => \GRLFPC2_0.N_1171\,
datae => \GRLFPC2_0.R.FSR.RD\(1),
datad => N_437,
datac => N_11,
datab => \GRLFPC2_0.N_3027\,
dataa => N_397);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_25_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30f0000020f00000")
port map (
combout => N_32903,
dataf => N_28634_1,
datae => N_34263_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_814\,
datac => N_32727_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A24_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0c0c0c0f0000000")
port map (
combout => N_32899,
dataf => N_33436_1,
datae => N_34341_1,
datad => N_28658_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A24_0\(55),
datab => N_32946);
\GRLFPC2_0_R_FSR_TEM_RNO_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"b888b888fccc3000")
port map (
combout => \GRLFPC2_0.R.FSR.TEM_1_0_0__G1\,
dataf => \GRLFPC2_0.N_1171\,
datae => \GRLFPC2_0.R.FSR.TEM\(0),
datad => N_429,
datac => N_11,
datab => \GRLFPC2_0.N_3027\,
dataa => N_389);
\GRLFPC2_0_R_FSR_TEM_RNO_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"b888b888fccc3000")
port map (
combout => \GRLFPC2_0.R.FSR.TEM_1_0_4__G1\,
dataf => \GRLFPC2_0.N_1171\,
datae => \GRLFPC2_0.R.FSR.TEM\(4),
datad => N_433,
datac => N_11,
datab => \GRLFPC2_0.N_3027\,
dataa => N_393);
\GRLFPC2_0_R_FSR_TEM_RNO_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"b888b888fccc3000")
port map (
combout => \GRLFPC2_0.R.FSR.TEM_1_0_3__G1\,
dataf => \GRLFPC2_0.N_1171\,
datae => \GRLFPC2_0.R.FSR.TEM\(3),
datad => N_432,
datac => N_11,
datab => \GRLFPC2_0.N_3027\,
dataa => N_392);
\GRLFPC2_0_R_FSR_TEM_RNO_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"b888b888fccc3000")
port map (
combout => \GRLFPC2_0.R.FSR.TEM_1_0_1__G1\,
dataf => \GRLFPC2_0.N_1171\,
datae => \GRLFPC2_0.R.FSR.TEM\(1),
datad => N_430,
datac => N_11,
datab => \GRLFPC2_0.N_3027\,
dataa => N_390);
\GRLFPC2_0_R_FSR_TEM_RNO_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"b888b888fccc3000")
port map (
combout => \GRLFPC2_0.R.FSR.TEM_1_0_2__G1\,
dataf => \GRLFPC2_0.N_1171\,
datae => \GRLFPC2_0.R.FSR.TEM\(2),
datad => N_431,
datac => N_11,
datab => \GRLFPC2_0.N_3027\,
dataa => N_391);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_10_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000c000000")
port map (
combout => N_33032,
dataf => N_29262_1,
datae => N_33507_1,
datad => N_32738_1_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0_O2_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fe505050ee000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8666\,
dataf => N_33735_1,
datae => N_28857_1,
datad => N_33138_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1659\,
datab => N_32818_I,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0faf0f0c0eac0c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_5\,
dataf => N_33794,
datae => N_33070_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1595\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9514\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_493\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A8_3_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"8080800000000000")
port map (
combout => N_28253,
dataf => N_28634_1,
datae => N_28658_1,
datad => N_28263,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_1_30_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33b300a000a000a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_30__G2_1\,
dataf => N_33735_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1586\,
datad => N_33798_I,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1222_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_COMB_RS1_1_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"eaff40ffea004000")
port map (
combout => \GRLFPC2_0.COMB.RS1_1\(4),
dataf => \GRLFPC2_0.R.A.RS1\(4),
datae => N_71,
datad => N_13,
datac => \GRLFPC2_0.RS1V_0_SQMUXA\,
datab => N_82,
dataa => \GRLFPC2_0.N_951\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_9_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cc005050dc50")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_8_1\,
dataf => N_34341_1,
datae => N_33178,
datad => N_29366_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_32_1\(58),
datab => N_33668_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff000fccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1028\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_473\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1586\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9600\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9511\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_15_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff02")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_15__G2_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9349\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8834\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9375\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_797\,
datab => N_33436_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11810_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffaeaa0c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_2__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19\(9),
datae => N_33794,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9502\,
datac => N_33140_1,
datab => N_28222_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1713\);
\GRLFPC2_0_COMB_RS1_1_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"eaff40ffea004000")
port map (
combout => \GRLFPC2_0.COMB.RS1_1\(3),
dataf => \GRLFPC2_0.R.A.RS1\(3),
datae => N_70,
datad => N_13,
datac => \GRLFPC2_0.RS1V_0_SQMUXA\,
datab => N_81,
dataa => \GRLFPC2_0.N_951\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A23_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0000000300000")
port map (
combout => N_33895,
dataf => N_32723_1,
datae => N_32858_1,
datad => N_28921_1,
datac => N_32791_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84));
\GRLFPC2_0_COMB_RS1_1_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"eaff40ffea004000")
port map (
combout => \GRLFPC2_0.COMB.RS1_1\(1),
dataf => \GRLFPC2_0.R.A.RS1\(1),
datae => N_68,
datad => N_13,
datac => \GRLFPC2_0.RS1V_0_SQMUXA\,
datab => N_79,
dataa => \GRLFPC2_0.N_951\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_0_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"88008a0000000a00")
port map (
combout => N_33022,
dataf => N_33507_1,
datae => N_33447_1,
datad => N_28560_2,
datac => N_33111,
datab => N_34195_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79));
\GRLFPC2_0_COMB_RS1_1_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"eaff40ffea004000")
port map (
combout => \GRLFPC2_0.COMB.RS1_1\(2),
dataf => \GRLFPC2_0.R.A.RS1\(2),
datae => N_69,
datad => N_13,
datac => \GRLFPC2_0.RS1V_0_SQMUXA\,
datab => N_80,
dataa => \GRLFPC2_0.N_951\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"dccccccc50000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_2\,
dataf => N_32738_1,
datae => N_33070_1,
datad => N_32782_1,
datac => N_28857_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1659\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffc0c0c0ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_719\,
datae => N_33652_1,
datad => N_32840_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1672\,
datab => N_28250_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_8_RNIK3437_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff75303030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1053\,
datae => N_34263_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1592\,
datac => N_32974_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_816\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000f444")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_758\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8556\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
datad => N_34341_1,
datac => N_33607_1,
datab => N_33718_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_6: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fddff72aa8dff77f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10864\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10879\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10878\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0_RNI9PIC_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff03")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_8__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9349\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9418\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_0\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_525\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_648\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff88ffffff80")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_12\,
dataf => N_33297_1,
datae => N_32732,
datad => N_32788,
datac => N_32796_3,
datab => N_32981_1,
dataa => N_33984_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_35_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000031300000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1492\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_429\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_I_O2_3_0\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_15_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f9f2fbf4fdf6ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(15),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(40),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_238_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0ff000eeeeeeee")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_238__G2_0_7736_I_0\,
dataf => \GRLFPC2_0.FPI.LDOP_0\,
datae => \GRLFPC2_0.FPI.OP2\(58),
datad => \GRLFPC2_0.FPI.OP2\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_40_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f2f4f6f9fbfdff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(40),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(16),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(15),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIA2RF_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0ff000eeeeeeee")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__G2_0_7550_I_0\,
dataf => \GRLFPC2_0.FPI.LDOP_0\,
datae => \GRLFPC2_0.FPI.OP2\(52),
datad => \GRLFPC2_0.FPI.OP2\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f2f9fbf4f6fdff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(13),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(42),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(43),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNI49VG_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0ff000eeeeeeee")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_243__G2_0_7581_I_0\,
dataf => \GRLFPC2_0.FPI.LDOP_0\,
datae => \GRLFPC2_0.FPI.OP2\(53),
datad => \GRLFPC2_0.FPI.OP2\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_237_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0ff000eeeeeeee")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_237__G2_0_7767_I_0\,
dataf => \GRLFPC2_0.FPI.LDOP_0\,
datae => \GRLFPC2_0.FPI.OP2\(59),
datad => \GRLFPC2_0.FPI.OP2\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_46_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f8f2faf5fdf7ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(46),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(10),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_239_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0ff000eeeeeeee")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_239__G2_0_7705_I_0\,
dataf => \GRLFPC2_0.FPI.LDOP_0\,
datae => \GRLFPC2_0.FPI.OP2\(57),
datad => \GRLFPC2_0.FPI.OP2\(60),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f9f2fbf4fdf6ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(10),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(45),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f2f4f6f9fbfdff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(42),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(14),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_16_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f2f4f6f9fbfdff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(16),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(40),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(39),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_14_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f2f9fbf4f6fdff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(14),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(41),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(43),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f4f8fcf3f7fbff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(49),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNI69VG_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0ff000eeeeeeee")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_241__G2_0_7643_I_0\,
dataf => \GRLFPC2_0.FPI.LDOP_0\,
datae => \GRLFPC2_0.FPI.OP2\(55),
datad => \GRLFPC2_0.FPI.OP2\(58),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f9f2fbf4fdf6ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(39),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(16),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_242_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0ff000eeeeeeee")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_242__G2_0_7612_I_0\,
dataf => \GRLFPC2_0.FPI.LDOP_0\,
datae => \GRLFPC2_0.FPI.OP2\(54),
datad => \GRLFPC2_0.FPI.OP2\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f9f4fdf2fbf6ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(17),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(40),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f8f2faf5fdf7ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(34),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(22),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(23),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(22),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f8f2faf5fdf7ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(18),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(38),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(39),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_R_E_STDATA_RNO_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"88f088ff88f08800")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_0__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(32),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.R.FSR.CEXC\(0),
datab => \GRLFPC2_0.R.I.INST\(0),
dataa => \GRLFPC2_0.N_91\);
\GRLFPC2_0_R_STATE_RNO_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000040c0000044cc")
port map (
combout => \GRLFPC2_0.R.STATE_0_0_0__G1\,
dataf => \GRLFPC2_0.N_1495\,
datae => \GRLFPC2_0.V.STATE_1_SQMUXA_3\,
datad => CPO_EXCZ,
datac => \GRLFPC2_0.R.STATE\(0),
datab => \GRLFPC2_0.N_1667\,
dataa => N_15);
\GRLFPC2_0_R_E_STDATA_RNO_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"88f088ff88f08800")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_1__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(33),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.R.FSR.CEXC\(1),
datab => \GRLFPC2_0.R.I.INST\(1),
dataa => \GRLFPC2_0.N_91\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_43_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f9f4fdf2fbf6ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(43),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(14),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(12),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_41_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f9f2fbf4fdf6ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(41),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(14),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(16),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0aaaaccccff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_ENA_67_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"060606060606ff00")
port map (
combout => N_38487,
dataf => \GRLFPC2_0.FPI.START\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(67),
datac => N_66,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7226\,
dataa => N_72);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_240_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0ff000eeeeeeee")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_240__G2_0_7674_I_0\,
dataf => \GRLFPC2_0.FPI.LDOP_0\,
datae => \GRLFPC2_0.FPI.OP2\(56),
datad => \GRLFPC2_0.FPI.OP2\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_5_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000a08000008080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1515\,
dataf => N_35132,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_492\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_429\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1637\,
datab => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_9_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"50d872fa55dd77ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(9),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(9),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_245_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"afaf00cca0a000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(245),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(12),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10530\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3639\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(245),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(232));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_0_0_TZ: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cc00cc00fff0ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_TZ\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1855\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_513\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_877_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_551\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_O2_0_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f400f400fffff555")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_402\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1855\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1730\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1566\,
datab => N_33652_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(66));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_250_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000fc30fc30")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(250),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10530\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10524\,
datad => \GRLFPC2_0.FPI.OP1\(62),
datac => \GRLFPC2_0.FPI.OP1\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_RNI217V_251_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000fc30fc30")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(251),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10530\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10523\,
datad => \GRLFPC2_0.FPI.OP1\(61),
datac => \GRLFPC2_0.FPI.OP1\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_RNI117V_252_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000fc30fc30")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(252),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10530\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10522\,
datad => \GRLFPC2_0.FPI.OP1\(60),
datac => \GRLFPC2_0.FPI.OP1\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_253_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000fc30fc30")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(253),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10530\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10521\,
datad => \GRLFPC2_0.FPI.OP1\(59),
datac => \GRLFPC2_0.FPI.OP1\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_254_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000fc30fc30")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(254),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10530\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10520\,
datad => \GRLFPC2_0.FPI.OP1\(58),
datac => \GRLFPC2_0.FPI.OP1\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_255_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000fc30fc30")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(255),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10530\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10519\,
datad => \GRLFPC2_0.FPI.OP1\(57),
datac => \GRLFPC2_0.FPI.OP1\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_RNI4T6V_256_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000fc30fc30")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(256),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10530\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10518\,
datad => \GRLFPC2_0.FPI.OP1\(56),
datac => \GRLFPC2_0.FPI.OP1\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_41_RNIJ4M71_257_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcc3300f0f0f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(257),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10530\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10503\,
datad => \GRLFPC2_0.FPO.EXP\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\(257),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26));
\GRLFPC2_0_R_E_STDATA_RNO_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0ccf0fff000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_2__G1\,
dataf => \GRLFPC2_0.R.A.AFSR\,
datae => \GRLFPC2_0.FPI.OP1\(34),
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_3052\,
datab => \GRLFPC2_0.R.FSR.CEXC\(2));
\GRLFPC2_0_R_E_STDATA_RNO_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3c0fffff3c00000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_3__G1\,
dataf => \GRLFPC2_0.N_3086\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.R.I.PC\(3),
datac => \GRLFPC2_0.R.I.INST\(3),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_R_E_STDATA_RNO_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0ccf0fff000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_4__G1\,
dataf => \GRLFPC2_0.R.A.AFSR\,
datae => \GRLFPC2_0.FPI.OP1\(36),
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_3054\,
datab => \GRLFPC2_0.R.FSR.CEXC\(4));
\GRLFPC2_0_R_E_STDATA_RNO_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0fff0ccf000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_5__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(37),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_3433\,
datab => \GRLFPC2_0.R.FSR.AEXC\(0));
\GRLFPC2_0_R_E_STDATA_RNO_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0fff0ccf000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_6__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(38),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_3056\,
datab => \GRLFPC2_0.R.FSR.AEXC\(1));
\GRLFPC2_0_R_E_STDATA_RNO_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3c0fffff3c00000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_7__G1\,
dataf => \GRLFPC2_0.N_3090\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.R.I.PC\(7),
datac => \GRLFPC2_0.R.I.INST\(7),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_R_E_STDATA_RNO_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3c0fffff3c00000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_8__G1\,
dataf => \GRLFPC2_0.N_3091\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.R.I.PC\(8),
datac => \GRLFPC2_0.R.I.INST\(8),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_R_E_STDATA_RNO_9_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0fff0ccf000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_9__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(41),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_3059\,
datab => \GRLFPC2_0.R.FSR.AEXC\(4));
\GRLFPC2_0_R_E_STDATA_RNO_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3c0fffff3c00000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_10__G1\,
dataf => \GRLFPC2_0.N_3093\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.R.I.PC\(10),
datac => \GRLFPC2_0.R.I.INST\(10),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_R_E_STDATA_RNO_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0fff0ccf000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_11__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(43),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_3434\,
datab => CPO_CCZ(1));
\GRLFPC2_0_R_E_STDATA_RNO_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000f0fff000f000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_12__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(44),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_3435\);
\GRLFPC2_0_R_E_STDATA_RNO_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ccffccf0cc00")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_13__G1\,
dataf => \GRLFPC2_0.N_71\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_76_I\,
datab => \GRLFPC2_0.N_3436\);
\GRLFPC2_0_R_E_STDATA_RNO_14_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3c0fffff3c00000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_14__G1\,
dataf => \GRLFPC2_0.N_3097\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.R.I.PC\(14),
datac => \GRLFPC2_0.R.I.INST\(14),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_R_E_STDATA_RNO_15_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000f0fff000f000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_15__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(47),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_3437\);
\GRLFPC2_0_R_E_STDATA_RNO_16_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3c0fffff3c00000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_16__G1\,
dataf => \GRLFPC2_0.N_3099\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.N_3423\,
datac => \GRLFPC2_0.R.I.INST\(16),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_R_E_STDATA_RNO_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0fff0fff0fff000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_17__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(49),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_3439\);
\GRLFPC2_0_R_E_STDATA_RNO_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3c0fffff3c00000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_18__G1\,
dataf => \GRLFPC2_0.N_3101\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.N_3425\,
datac => \GRLFPC2_0.R.I.INST\(18),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_R_E_STDATA_RNO_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000f0fff000f000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_19__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(51),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_3069\);
\GRLFPC2_0_R_E_STDATA_RNO_20_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3c0fffff3c00000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_20__G1\,
dataf => \GRLFPC2_0.N_3103\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.N_3426\,
datac => \GRLFPC2_0.R.I.INST\(20),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_R_E_STDATA_RNO_21_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000f0fff000f000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_21__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(53),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_3442\);
\GRLFPC2_0_R_E_STDATA_RNO_22_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0fff0ccf000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_22__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(54),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_3443\,
datab => \GRLFPC2_0.R.FSR.NONSTD\);
\GRLFPC2_0_R_E_STDATA_RNO_23_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3c0fffff3c00000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_23__G1\,
dataf => \GRLFPC2_0.N_3106\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.N_3429\,
datac => \GRLFPC2_0.R.I.INST\(23),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_R_E_STDATA_RNO_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0fff0ccf000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_24__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(56),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_3445\,
datab => \GRLFPC2_0.R.FSR.TEM\(1));
\GRLFPC2_0_R_E_STDATA_RNO_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3c0fffff3c00000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_25__G1\,
dataf => \GRLFPC2_0.N_3108\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.R.I.PC\(25),
datac => \GRLFPC2_0.R.I.INST\(25),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_R_E_STDATA_RNO_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3c0fffff3c00000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_26__G1\,
dataf => \GRLFPC2_0.N_3109\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.R.I.PC\(26),
datac => \GRLFPC2_0.R.I.INST\(26),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_R_E_STDATA_RNO_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0fff0ccf000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_27__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(59),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_3077\,
datab => \GRLFPC2_0.R.FSR.TEM\(4));
\GRLFPC2_0_R_E_STDATA_RNO_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000f0fff000f000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_28__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(60),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_3078\);
\GRLFPC2_0_R_E_STDATA_RNO_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000f0fff000f000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_29__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(61),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_3079\);
\GRLFPC2_0_R_E_STDATA_RNO_30_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccf0fff0ccf000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_30__G1\,
dataf => \GRLFPC2_0.FPI.OP1\(62),
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.A.AFQ\,
datac => \GRLFPC2_0.N_3446\,
datab => \GRLFPC2_0.R.FSR.RD\(0));
\GRLFPC2_0_R_E_STDATA_RNO_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3c0fffff3c00000")
port map (
combout => \GRLFPC2_0.R.E.STDATA_1_0_31__G1\,
dataf => \GRLFPC2_0.N_3114\,
datae => \GRLFPC2_0.R.A.AFQ\,
datad => \GRLFPC2_0.N_3432\,
datac => \GRLFPC2_0.R.I.INST\(31),
datab => \GRLFPC2_0.N_91\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_27_S: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(49));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_BUSYMULXFF_UN2_TEMP_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.BUSYMULXFF.UN2_TEMP_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(68),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(70));
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_0_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfcfcfcfcfc0cfcf")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV_0\(4),
dataf => \GRLFPC2_0.N_1133\,
datae => \GRLFPC2_0.N_1171\,
datad => N_375,
datac => \GRLFPC2_0.N_1517\,
datab => N_415);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cc00fc00cc00ff00")
port map (
combout => \GRLFPC2_0.R.FSR.AEXC_1_0_4__I0_I_0\,
dataf => \GRLFPC2_0.V.FSR.CEXC_0_SQMUXA\,
datae => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA\,
datad => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV_0\(4),
datac => \GRLFPC2_0.R.I.EXC\(4),
datab => \GRLFPC2_0.R.FSR.AEXC\(4));
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c0f0ccff00000000")
port map (
combout => \GRLFPC2_0.R.FSR.CEXC_1_0_0__I0_I_1\,
dataf => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_1\(0),
datae => \GRLFPC2_0.V.FSR.CEXC_0_SQMUXA\,
datad => \GRLFPC2_0.V.FSR.CEXC_3_SQMUXA\,
datac => \GRLFPC2_0.R.I.EXC\(0),
datab => \GRLFPC2_0.R.FSR.CEXC\(0));
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c0f0ccff00000000")
port map (
combout => \GRLFPC2_0.R.FSR.CEXC_1_0_1__I0_I_0\,
dataf => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_1\(1),
datae => \GRLFPC2_0.V.FSR.CEXC_0_SQMUXA\,
datad => \GRLFPC2_0.V.FSR.CEXC_3_SQMUXA\,
datac => \GRLFPC2_0.R.I.EXC\(1),
datab => \GRLFPC2_0.R.FSR.CEXC\(1));
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c0f0ccff00000000")
port map (
combout => \GRLFPC2_0.R.FSR.CEXC_1_0_3__I0_I_0\,
dataf => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_1\(3),
datae => \GRLFPC2_0.V.FSR.CEXC_0_SQMUXA\,
datad => \GRLFPC2_0.V.FSR.CEXC_3_SQMUXA\,
datac => \GRLFPC2_0.R.I.EXC\(3),
datab => \GRLFPC2_0.R.FSR.CEXC\(3));
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c0f0ccff00000000")
port map (
combout => \GRLFPC2_0.R.FSR.CEXC_1_0_4__I0_I_1\,
dataf => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_1\(4),
datae => \GRLFPC2_0.V.FSR.CEXC_0_SQMUXA\,
datad => \GRLFPC2_0.V.FSR.CEXC_3_SQMUXA\,
datac => \GRLFPC2_0.R.I.EXC\(4),
datab => \GRLFPC2_0.R.FSR.CEXC\(4));
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_0_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfcfcfcfcfc0cfcf")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV_0\(0),
dataf => \GRLFPC2_0.N_1133\,
datae => \GRLFPC2_0.N_1171\,
datad => N_371,
datac => \GRLFPC2_0.N_1517\,
datab => N_411);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cc00fc00cc00ff00")
port map (
combout => \GRLFPC2_0.R.FSR.AEXC_1_0_0__I0_I_0\,
dataf => \GRLFPC2_0.V.FSR.CEXC_0_SQMUXA\,
datae => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA\,
datad => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV_0\(0),
datac => \GRLFPC2_0.R.I.EXC\(0),
datab => \GRLFPC2_0.R.FSR.AEXC\(0));
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_0_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfcfcfcfcfc0cfcf")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV_0\(2),
dataf => \GRLFPC2_0.N_1133\,
datae => \GRLFPC2_0.N_1171\,
datad => N_373,
datac => \GRLFPC2_0.N_1517\,
datab => N_413);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cc00fc00cc00ff00")
port map (
combout => \GRLFPC2_0.R.FSR.AEXC_1_0_2__I0_I_0\,
dataf => \GRLFPC2_0.V.FSR.CEXC_0_SQMUXA\,
datae => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA\,
datad => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV_0\(2),
datac => \GRLFPC2_0.R.I.EXC\(2),
datab => \GRLFPC2_0.R.FSR.AEXC\(2));
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_0_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfcfcfcfcfc0cfcf")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV_0\(3),
dataf => \GRLFPC2_0.N_1133\,
datae => \GRLFPC2_0.N_1171\,
datad => N_374,
datac => \GRLFPC2_0.N_1517\,
datab => N_414);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cc00fc00cc00ff00")
port map (
combout => \GRLFPC2_0.R.FSR.AEXC_1_0_3__I0_I_1\,
dataf => \GRLFPC2_0.V.FSR.CEXC_0_SQMUXA\,
datae => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA\,
datad => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV_0\(3),
datac => \GRLFPC2_0.R.I.EXC\(3),
datab => \GRLFPC2_0.R.FSR.AEXC\(3));
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_0_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfcfcfcfcfc0cfcf")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV_0\(1),
dataf => \GRLFPC2_0.N_1133\,
datae => \GRLFPC2_0.N_1171\,
datad => N_372,
datac => \GRLFPC2_0.N_1517\,
datab => N_412);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cc00fc00cc00ff00")
port map (
combout => \GRLFPC2_0.R.FSR.AEXC_1_0_1__I0_I_1\,
dataf => \GRLFPC2_0.V.FSR.CEXC_0_SQMUXA\,
datae => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA\,
datad => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV_0\(1),
datac => \GRLFPC2_0.R.I.EXC\(1),
datab => \GRLFPC2_0.R.FSR.AEXC\(1));
GRLFPC2_0_V_STATE_0_SQMUXA_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000000000")
port map (
combout => \GRLFPC2_0.N_1517\,
dataf => N_398,
datae => N_399,
datad => N_400);
GRLFPC2_0_COMB_ANNULFPU_1_U_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffc30")
port map (
combout => \GRLFPC2_0.COMB.ANNULFPU_1\,
dataf => \GRLFPC2_0.COMB.ANNULFPU_1_U_0_0\,
datae => \GRLFPC2_0.N_3491\,
datad => \GRLFPC2_0.R.X.FPOP\,
datac => \GRLFPC2_0.R.X.SEQERR\,
datab => \GRLFPC2_0.N_1105\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_7_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0f000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_403\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_A2_7_1\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856\,
datac => N_59);
GRLFPC2_0_COMB_V_A_AFSR_1_0_A2_1_0_RNIM8CH1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => \GRLFPC2_0.R.A.AFSR\,
dataf => \GRLFPC2_0.N_552_1_0\,
datae => \GRLFPC2_0.R.E.AFQ_RET_0_0_G1_5\,
datad => \GRLFPC2_0.FPCI_O\(59),
datac => \GRLFPC2_0.FPCI_O\(62),
datab => \GRLFPC2_0.FPCI_O\(58));
\GRLFPC2_0_R_A_AFQ_RET_RNIIOHR_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000f000000")
port map (
combout => \GRLFPC2_0.R.E.AFQ_RET_0_0_G1_3\,
dataf => \GRLFPC2_0.FPCI_O\(58),
datae => \GRLFPC2_0.FPCI_O\(60),
datad => \GRLFPC2_0.FPCI_O\(63),
datac => \GRLFPC2_0.FPCI_O\(61));
\GRLFPC2_0_R_A_AFQ_RET_RNID06U2_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000000000000000")
port map (
combout => \GRLFPC2_0.R.A.AFQ\,
dataf => \GRLFPC2_0.R.E.AFQ_RET_0_0_G1_5\,
datae => \GRLFPC2_0.N_202\,
datad => \GRLFPC2_0.R.E.AFQ_RET_0_0_G1_3\,
datac => \GRLFPC2_0.FPCI_O\(59),
datab => \GRLFPC2_0.FPCI_O\(62));
GRLFPC2_0_COMB_V_A_AFSR_1_0_A2_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff0000000000")
port map (
combout => \GRLFPC2_0.N_552_1_0\,
dataf => \GRLFPC2_0.N_202\,
datae => \GRLFPC2_0.FPCI_O\(61),
datad => \GRLFPC2_0.FPCI_O\(63));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIOCHD_64_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW_2\(65),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3926\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(68),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(64));
\GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c0f0ccff00000000")
port map (
combout => \GRLFPC2_0.R.FSR.CEXC_1_0_2__I0_I_1\,
dataf => \GRLFPC2_0.COMB.V.FSR.CEXC_1_IV_1\(2),
datae => \GRLFPC2_0.V.FSR.CEXC_0_SQMUXA\,
datad => \GRLFPC2_0.V.FSR.CEXC_3_SQMUXA\,
datac => \GRLFPC2_0.R.I.EXC\(2),
datab => \GRLFPC2_0.R.FSR.CEXC\(2));
GRLFPC2_0_R_I_EXEC_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f30000ffff0000")
port map (
combout => N_37428,
dataf => N_37318_1,
datae => \GRLFPC2_0.R.I.EXEC_0_0_G1_0_7945_I_3\,
datad => \GRLFPC2_0.COMB.ISFPOP2_1\,
datac => \GRLFPC2_0.R.X.LD\,
datab => \GRLFPC2_0.R.I.V\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_2_RNITA48_0_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0f33f0f0f0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(374),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(0));
\GRLFPC2_0_R_I_EXC_RNO_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f0000000000000")
port map (
combout => \GRLFPC2_0.R.I.EXC_2_0_2__G2\,
dataf => \GRLFPC2_0.R.I.EXC_MB\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(40),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(38));
\GRLFPC2_0_R_A_RF2REN_RNO_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000fff00000")
port map (
combout => N_37432,
dataf => N_37387,
datae => \GRLFPC2_0.N_951\,
datad => \GRLFPC2_0.N_77_1\,
datac => N_53);
GRLFPC2_0_R_MK_BUSY_RET_4_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000c000000000")
port map (
combout => \GRLFPC2_0.N_2111\,
dataf => \GRLFPC2_0.R.MK.RST_4\,
datae => \GRLFPC2_0.R.MK.RST2\,
datad => \GRLFPC2_0.R.MK.RST2_O\,
datac => \GRLFPC2_0.COMB.ANNULFPU_1_O\,
datab => N_11);
GRLFPC2_0_R_MK_BUSY2_RET_1_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ff00")
port map (
combout => \GRLFPC2_0.N_2105\,
dataf => \GRLFPC2_0.N_3545\,
datae => \GRLFPC2_0.COMB.ANNULFPU_1_O_0\,
datad => N_11);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_10_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff000000f0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1520\,
dataf => N_35132,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1637\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1771\,
datac => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_8_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1518\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1493\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1492\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_451\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_492\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_6_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cc000000c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1516\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1836\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_492\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1636\,
datac => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_1_A2_7_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_A2_1_A2_7\(83),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1518\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_A2_1_A2_2\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1516\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1519\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_1_A2_9_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000007f00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_A2_1_A2_9\(83),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_A2_1_A2_7\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1515\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1520\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1844\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1636\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1771\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_7_0_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc300000fc30fc30")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_A2_7_0\(83),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_A2_7_8923_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_492\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_504\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_7_2_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff00cf00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_A2_7_2\(83),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1505\,
datae => N_35132,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_A2_7_0\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1637\,
datab => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_41_0_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0ffff03f3ffff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_A2_41_0\(83),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_I_O2_3_0\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_41_2_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_A2_41_2\(83),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_451\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_A2_41_0\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1677\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1770\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_41_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000003f000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1505\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1495\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_A2_41_2\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233));
GRLFPC2_0_RS2_0_SQMUXA_0_0_A2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000000000")
port map (
combout => \GRLFPC2_0.N_951\,
dataf => \GRLFPC2_0.N_3462\,
datae => N_76,
datad => N_74,
datac => N_83,
datab => N_73);
GRLFPC2_0_R_A_RDD_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f0000000000000")
port map (
combout => \GRLFPC2_0.R.A.RDD_0_0_G1\,
dataf => \GRLFPC2_0.COMB.RDD_1.N_12\,
datae => N_77,
datad => N_75,
datac => N_84);
GRLFPC2_0_COMB_LOCK_1_I: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000030000")
port map (
combout => CPO_LDLOCKZ,
dataf => \GRLFPC2_0.R.STATE\(1),
datae => \GRLFPC2_0.N_3477_1_I\,
datad => N_88,
datac => \GRLFPC2_0.R.STATE\(0),
datab => N_87);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_19_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fcf000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_19\(60),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_3\(60),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_4\(60),
datad => N_33146_1,
datac => N_33718_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_8_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcffffffffcfffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_8\(60),
dataf => N_33144_1,
datae => N_28250_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_2_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000003fffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_2\(60),
dataf => N_33729,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_531\,
datad => N_33721_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"2000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__I0_I_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_18\(60),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_20\(60),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_19\(60),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_17\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9166\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_16\(60));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_17_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_17\(11),
dataf => N_33968,
datae => N_33973,
datad => N_33971,
datac => N_33976,
datab => N_33974);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_0_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000003fffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_0\(11),
dataf => N_33967,
datae => N_33436_1,
datad => N_33899_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_16_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000030000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_16\(11),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_0\(11),
datae => N_33987,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_3\(11),
datac => N_33975,
datab => N_33982);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_11_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000003fff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_11\(11),
dataf => N_33966,
datae => N_33970,
datad => N_28492_1,
datac => N_33988_4,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_21_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"4000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_21\(11),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_11\(11),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_6\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_13\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_7\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_12\(11),
dataa => N_33972);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fc00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_11__I0_I_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_21\(11),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_17\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_16\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_525\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_648\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_11_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00003fff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_11\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_2\(47),
datae => N_33733,
datad => N_32844_2,
datac => N_33436_1,
datab => N_33138_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_8_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f3ffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_8\(47),
dataf => N_34255,
datae => N_32844_2,
datad => N_32796_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_7_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff3fff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_7\(47),
dataf => N_34259,
datae => N_33436_1,
datad => N_32858_1,
datac => N_28549_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_14_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3fff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_14\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_7\(47),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_0\(47),
datad => N_34272_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_20_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_20\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_14\(47),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_8\(47),
datad => N_32844_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_10_TZ\(47),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_1_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"033333330fffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_1\(47),
dataf => N_33436_1,
datae => N_33138_1,
datad => N_32786_1,
datac => N_28261_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_15_0\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_18_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000333")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_18\(47),
dataf => N_32981,
datae => N_34260,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_8_0\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_8_1\(47),
datab => N_34268);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_22_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000030000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_22\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_18\(47),
datae => N_34271,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_1\(47),
datac => N_34262,
datab => N_34279);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_48__I0_I_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_20\(47),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_22\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_11\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_9\(47),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1135\,
dataa => N_34254);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN2_NOTDECODEDUNIMP: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccfffcffccffccff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3926\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_475\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(66),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(67),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(64));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A26_1_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0033003000000000")
port map (
combout => N_33966,
dataf => N_29653_1,
datae => N_32979_1,
datad => N_28250_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A26_2_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000c000f03")
port map (
combout => N_33967,
dataf => N_33055,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A26_6_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000003000000")
port map (
combout => N_33971,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_719\,
datae => N_34239_I,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A26_8_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000c0000000c000")
port map (
combout => N_33973,
dataf => N_33436_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_531\,
datad => N_33501_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A26_9_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => N_33974,
dataf => N_33652_1,
datae => N_32959_I,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_5_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000c000")
port map (
combout => N_34260,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_782\,
datae => N_33574_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_7_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => N_34262,
dataf => N_28264_1,
datae => N_34233,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_15_0_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_15_0\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A28_14_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000003000")
port map (
combout => N_33733,
dataf => N_34029,
datae => N_34239_I,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A8_5_0_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A8_5_0\(62),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A8_1_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0c0c0c000000000")
port map (
combout => N_28251,
dataf => N_32844_2,
datae => N_32982_1,
datad => N_28266_2,
datac => N_28251_1,
datab => N_28267);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_63_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff0fcf0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_2\,
dataf => N_28251,
datae => N_29653_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_797\,
datac => N_28252,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A8_5_0\(62));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffc0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_2\,
dataf => N_28210,
datae => N_33659_1,
datad => N_33436_1,
datac => N_28560_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A11_6_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"300c000000000000")
port map (
combout => N_28212,
dataf => N_29195_1,
datae => N_28212_1_0,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_0\,
datac => N_28212,
datab => N_28206,
dataa => N_28207);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000ccc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_531\,
datad => N_28226,
datac => N_28227,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_1_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000003cf00000000")
port map (
combout => N_33897,
dataf => N_33870,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_19\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_13\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_11\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_12\,
datac => N_33913,
datab => N_33912,
dataa => N_33900);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_10_0_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_10_0\(59),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_15\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_9\,
datae => N_33896,
datad => N_32727_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_2_1\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_12_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0330000000000000")
port map (
combout => N_33908,
dataf => N_32730_1,
datae => N_28921_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff40")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_19\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_15\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_7\,
datac => N_33735_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_5_1\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_37_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"030c000000000000")
port map (
combout => N_33654,
dataf => N_33436_1,
datae => N_33503_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A29_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3330000030300000")
port map (
combout => N_33643,
dataf => N_28266_2,
datae => N_28212_1,
datad => N_29366_1,
datac => N_33683,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_29_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3300300000000000")
port map (
combout => N_33646,
dataf => N_33735_1,
datae => N_33447_1,
datad => N_33503_1,
datac => N_33734_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_49_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => N_33666,
dataf => N_32982_1,
datae => N_33503_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_30_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000300000")
port map (
combout => N_33647,
dataf => N_28634_1,
datae => N_32982_1,
datad => N_33507_1,
datac => N_28261_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_20\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_22\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_13\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_12\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9397\,
dataa => N_33644);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_18_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_5\,
datad => N_33148,
datac => N_33130,
datab => N_33134);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A32_25_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => N_33149,
dataf => N_33659_1,
datae => N_32796_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_10_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000300000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_782\,
datae => N_32909_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_21\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_18_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_20\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_14\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_23\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_13_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_2_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0ccc0000000000")
port map (
combout => N_33210,
dataf => N_32979_1,
datae => N_33179,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00000c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_2\,
dataf => N_33229,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_719\,
datad => N_32727_1,
datac => N_32821,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_9_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000003c")
port map (
combout => N_33217,
dataf => N_33055,
datae => N_33004,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff00c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_9\,
dataf => N_33217,
datae => N_33224,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_719\,
datac => N_32796_2,
datab => N_28250_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_7_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000c300000000")
port map (
combout => N_33215,
dataf => N_32844_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_719\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_1_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000000030000000")
port map (
combout => N_33209,
dataf => N_32979_1,
datae => N_28222_1,
datad => N_32727_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_9_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffc0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_7\,
dataf => N_33209,
datae => N_33659_1,
datad => N_33436_1,
datac => N_28560_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_A28_11_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000ccf0000")
port map (
combout => N_33219,
dataf => N_33178,
datae => N_33253,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_10_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00c0ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_14\,
dataf => N_29653_1,
datae => N_33207,
datad => N_33503_1,
datac => N_33253,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_11_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00000030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_4\,
dataf => N_33208,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_782\,
datad => N_32818_I,
datac => N_28652_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_18\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_11\,
datad => N_33222_2,
datac => N_33179,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_22\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_18\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_13\,
datad => N_28658_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_16_TZ\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_22\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_16_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_20\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_9\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_36_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30c0000000000000")
port map (
combout => N_32914,
dataf => N_32738_1,
datae => N_32727_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_31_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c300000000000000")
port map (
combout => N_32909,
dataf => N_33436_1,
datae => N_34329_1,
datad => N_32909_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00c00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_2\,
dataf => N_32909,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_0_1\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffcfff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_12\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_10_TZ\,
datad => N_32902,
datac => N_32912,
datab => N_32946);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f3f000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_6\,
dataf => N_32979_1,
datae => N_33138_1,
datad => N_33607_1,
datac => N_33111,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_28_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0003000000000000")
port map (
combout => N_32906,
dataf => N_32844_2,
datae => N_34341_1,
datad => N_33368_1,
datac => N_32738_1_0,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_15\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_6\,
datad => N_32903,
datac => N_32906,
datab => N_33913);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_37_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000c30000")
port map (
combout => N_32915,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11641\,
datae => N_33607_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_17\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_15\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_12\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_9\,
datab => N_32921);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_9\,
dataf => N_34120,
datae => N_34117,
datad => N_32738_1,
datac => N_32723_1,
datab => N_34132_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_1_1_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"003f000c00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_1_1\(54),
dataf => N_32858_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff00c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_14\,
dataf => N_34123,
datae => N_34121,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11641\,
datac => N_29195_1,
datab => N_34133_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_2_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000300000000000")
port map (
combout => N_34113,
dataf => N_32738_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_719\,
datad => N_32723_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffc0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_4\,
dataf => N_34118,
datae => N_32723_1,
datad => N_32858_1,
datac => N_28250_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_19\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_18\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_15\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_7\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_9\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_17\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_19_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030000000000000")
port map (
combout => N_33847,
dataf => N_33543,
datae => N_33984_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_0_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000ccc0000")
port map (
combout => N_33828,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_797\,
datae => N_33543,
datad => N_33178,
datac => N_33111,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_5_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => N_33833,
dataf => N_29653_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_719\,
datad => N_34341_1,
datac => N_33111,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_11_0\,
dataf => N_33833,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_5\,
datad => N_33543,
datac => N_33838_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_15\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_11_0\,
datae => N_33828,
datad => N_33847,
datac => N_32904_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_11_TZ\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_7_1_0_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000c0c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_7_1\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_6_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000c00c0000")
port map (
combout => N_33834,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_531\,
datae => N_28227_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff000000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_1\,
dataf => N_33839,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_719\,
datad => N_33798_I,
datac => N_32980_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff8")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_15\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_13\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_10\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1374\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_1_0\(53),
dataa => N_33813);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_2_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c0c00000c0000000")
port map (
combout => N_33501,
dataf => N_33144_1,
datae => N_33501_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_14\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_0\,
datae => N_33518,
datad => N_33505,
datac => N_33501,
datab => N_33498);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_4_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"030f000000000000")
port map (
combout => N_33503,
dataf => N_33725_1,
datae => N_33503_1,
datad => N_33263_I,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_3_0_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_3_0\(52),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_5_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030003f00000000")
port map (
combout => N_33504,
dataf => N_28549_1,
datae => N_33263_I,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_604\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff000c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_10\,
dataf => N_33506,
datae => N_32730_1,
datad => N_33111,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_0_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000c00f000")
port map (
combout => N_33499,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datae => N_33725_1,
datad => N_32727_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffc0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_2\,
dataf => N_33499,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datad => N_28271_1,
datac => N_33507_1,
datab => N_28250_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_18\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_14\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8941\,
datab => N_33513,
dataa => N_33510);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff8")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_16\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_9\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_6\,
datad => N_34334,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_11\,
datab => N_34325_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0_1\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_16\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_11_0\,
dataa => N_34337);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff03000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1187\,
datae => N_32723_1,
datad => N_33146_1,
datac => N_32722_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_4\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_5\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_11\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1233\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1237\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1236\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff0c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_10\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_659\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1682\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_525\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9547\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_10\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_11\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_9\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_584\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1235\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1234\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_5_0_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f0000f0ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_5_0\(48),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_3_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000303300000000")
port map (
combout => N_34184,
dataf => N_33659_1,
datae => N_33548,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_531\,
datac => N_28658_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_7\,
dataf => N_34184,
datae => N_34182,
datad => N_33146_1,
datac => N_28564_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_5_0\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_2_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"003c000000000000")
port map (
combout => N_34183,
dataf => N_32844_3,
datae => N_33899_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_9_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000c0000000")
port map (
combout => N_34190,
dataf => N_32861_1,
datae => N_29071_1,
datad => N_32730_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_6_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c300000000000000")
port map (
combout => N_34187,
dataf => N_32861_1,
datae => N_28211_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_10\,
dataf => N_34180,
datae => N_34190,
datad => N_34187);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_18\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_10\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1053\,
datad => N_34191,
datac => N_34337,
datab => N_34195);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_18\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_13\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_14\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_6\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_948\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_5\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff0fc00cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_47__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1031\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9486\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_797\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9502\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1659\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_45_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c3c300000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2_1\,
dataf => N_32844_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9600\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9547\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_15_I_O2_RNI0MGR1_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f000fcccf000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9486\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_473\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_648\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_RNI0I772_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_758\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1194\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1758\,
datab => N_32974_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_6_0_A2_RNIC05N4_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f030c0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2_0\,
dataf => N_33070_1,
datae => N_32840_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9570\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_1_A2_RNI0MO35_41_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9166\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9165\,
datac => N_33794,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9486\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_41_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffccfc00f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_41__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1278\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9502\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_571\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9492\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9490\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_40_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff03")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_40__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_693\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_0_0\(39),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1744\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_571\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_814\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_0_0_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000cf03cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_0_0\(39),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9525\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0_1\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_39__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_39__G2_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_756\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_0_0\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1744\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_756\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1588\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1133\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_5_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cc3f000000000000")
port map (
combout => N_32727,
dataf => N_32727_1,
datae => N_32796_3,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_2_0_0_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_2_0_0\(36),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffc000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_9\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_4\,
datae => N_32722_1,
datad => N_32722_2,
datac => N_28730_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_13\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_9\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_3\,
datac => N_32729,
datab => N_32735);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_13\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_7\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9157\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_6\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_907\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_12\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_35_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c00c000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9198\,
dataf => N_34263_2,
datae => N_33123_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0fcf0ff00cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9525\,
datae => N_34341_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9502\,
datac => N_28658_1,
datab => N_32732_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff00c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1206\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1201\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\,
datac => N_28857_1,
datab => N_28564_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffcf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_11\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9418\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1586\,
datac => N_32732,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1757\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_11\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_769\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_9\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_5\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0c000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_2\,
dataf => N_32787,
datae => N_29653_1,
datad => N_33055,
datac => N_29518_1,
datab => N_32980_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000fccc0000cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_1\,
dataf => N_33340_I,
datae => N_33004,
datad => N_28564_2,
datac => N_32786_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A24_4_1\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00003000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datad => N_28857_1,
datac => N_33984_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_17\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_2\,
datad => N_32798,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1222_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_5_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000c0000000000")
port map (
combout => N_32783,
dataf => N_33507_1,
datae => N_28564_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_2_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000300030000")
port map (
combout => N_32780,
dataf => N_32861_1,
datae => N_32844_3,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff000000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_4\,
dataf => N_32780,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datad => N_32762_I,
datac => N_33984_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_16\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_4\,
datae => N_32785,
datad => N_32777,
datac => N_32783,
datab => N_32788);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_17\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_16\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_15\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9157\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1206\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_5_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cc000000c000")
port map (
combout => N_33289,
dataf => N_33074_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_531\,
datad => N_34254_1,
datac => N_28261_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_5_RNISF3Q8_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff30000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_2\,
dataf => N_33289,
datae => N_34340_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_7_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000f300")
port map (
combout => N_33291,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\,
datae => N_33548,
datad => N_32738_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_2_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000330000003000")
port map (
combout => N_33286,
dataf => N_32861_1,
datae => N_33548,
datad => N_33503_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_3_1_RNI6RFL8_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffff00ffc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_9\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_4\,
datae => N_33548,
datad => N_33590,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_3_1\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A17_RNI5JE79_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffec")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_11\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_9\,
datae => N_33297,
datad => N_33288,
datac => N_32861_1,
datab => N_33283,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_11_0\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_7_RNIH66B41_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_11\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_6\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_7\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_907\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A14_2_2_RNI5V397_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f0000c00fc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_17\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_525\,
datae => N_32840_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_7_RNIT7A53_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0300ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_6\,
dataf => N_28271_1,
datae => N_33578,
datad => N_28564_2,
datac => N_32727_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_5_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30fc000000000000")
port map (
combout => N_33576,
dataf => N_32844_2,
datae => N_28212_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_10_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000000000000000")
port map (
combout => N_33581,
dataf => N_32861_1,
datae => N_33548,
datad => N_33503_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_37_1_RNIP4K1Q_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_18\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_12\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_7\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_6\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_17\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_0_30_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000f000f000fccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_30__G2_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_525\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9509\,
datac => N_33369_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_1_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1388\,
datae => N_33589,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1389\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9503\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9509\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_0_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1832\,
datad => N_32782_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1592\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_30_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffcccfffff000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_759\,
dataf => N_34271,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_907\,
datad => N_33794,
datac => N_34040_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cf0fcc00cc00cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_0\,
dataf => N_32979_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9517\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_8_0\(47),
datac => N_33263_I,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_8_1\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_17_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000003000000000")
port map (
combout => N_33588,
dataf => N_29071_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_23_0_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f000000330000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_23_0\(27),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_29_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0330000000000000")
port map (
combout => N_33358,
dataf => N_33074_1,
datae => N_33368_1,
datad => N_33144_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_28_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000003c00000000")
port map (
combout => N_33357,
dataf => N_32844_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_719\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_33_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000030f")
port map (
combout => N_33362,
dataf => N_33548,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_797\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_26_0_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00000000ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_26_0\(27),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffc0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_1\,
dataf => N_33362,
datae => N_33144_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_26_0\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_17\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_5\,
datac => N_33357,
datab => N_33358,
dataa => N_33351);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff000000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_4\,
dataf => N_33360,
datae => N_32844_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_719\,
datac => N_28658_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffcf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_19\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_13\,
datad => N_33794,
datac => N_33369,
datab => N_28222_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_17\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_19\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_10\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_9\,
datab => N_33373,
dataa => N_33359);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffc0c0c0c0c0c0c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_2\,
dataf => N_32738_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9525\,
datad => N_28266_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9600\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11810_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_8\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_584\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1038\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_24__G2_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8666\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9327\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_525\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_816\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_24__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_24__G2_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9608\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9665\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9645\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9607\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_21_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffcccf000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_21__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9158\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9486\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9525\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9498\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9492\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_26_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f0000000c00000")
port map (
combout => N_33428,
dataf => N_32730_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1607\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_23_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f030000000000000")
port map (
combout => N_33425,
dataf => N_32738_1,
datae => N_33140_1,
datad => N_32786_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_28_0_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff0000000000ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_28_0\(19),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_28_0_RNIH5OU2_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccc0cc00c0c00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_0\,
dataf => N_32738_1,
datae => N_29366_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_28_0\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datab => N_28730_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_32_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000c000000")
port map (
combout => N_33434,
dataf => N_33543,
datae => N_34254_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_37_0_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_37_0\(19),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_34_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => N_33436,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_782\,
datae => N_33436_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_37_0_RNIVQ6D6_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00003000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_6\,
dataf => N_33436,
datae => N_33146_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_37_0\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_38_RNIS7TU1_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffc0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_5\,
dataf => N_33440,
datae => N_28264_1,
datad => N_33574_1,
datac => N_33146_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_25_RNI6U5R8_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_18\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_5\,
datad => N_33427,
datac => N_33434,
datab => N_33444);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_33_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000033300000000")
port map (
combout => N_33435,
dataf => N_28264_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_31_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c030000000000000")
port map (
combout => N_33433,
dataf => N_33507_1,
datae => N_32722_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_27_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000f0")
port map (
combout => N_33429,
dataf => N_33411,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_35_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0003000000000000")
port map (
combout => N_33437,
dataf => N_33543,
datae => N_32723_1,
datad => N_33081_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_24_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000c000000")
port map (
combout => N_33426,
dataf => N_32738_1,
datae => N_33507_1,
datad => N_33140_1,
datac => N_33368_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_24_RNI415I_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff000c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_10\,
dataf => N_33426,
datae => N_33437,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\,
datac => N_33138_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_15_1\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_30_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0c00000c000000")
port map (
combout => N_33432,
dataf => N_33368_1,
datae => N_28564_2,
datad => N_33503_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_27_RNI5OHIA_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_20\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_10\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_9\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_3\,
datac => N_33447,
datab => N_33435,
dataa => N_33429);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_23_RNI2JCVR_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_20\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_18\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_8\,
datac => N_33431,
datab => N_33425,
dataa => N_33428);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_2_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000003000000000")
port map (
combout => N_33069,
dataf => N_33055,
datae => N_33004,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00003000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_10\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_6\,
datae => N_32723_1,
datad => N_33146_1,
datac => N_33061,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_1_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3033000000000000")
port map (
combout => N_33068,
dataf => N_33436_1,
datae => N_32858_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_3_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00003f0000000000")
port map (
combout => N_33070,
dataf => N_33070_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\,
datad => N_32723_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_7\,
dataf => N_33070,
datae => N_33073,
datad => N_33071,
datac => N_28857_1,
datab => N_33138_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_11\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_7\,
datae => N_33076,
datad => N_32723_1,
datac => N_33140_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9492\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_10\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_11\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1304\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_9_RNIEEKN_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_12\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9397\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_544\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1054\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1586\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9492\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_RNI24HLF_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff03")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_10\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_6\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9368\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_525\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_814\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_10\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_12\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8714\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9349\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9373\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_RNIHQCC5_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_16__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_693\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_16__G2_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_571\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8619\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_15_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff0c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_15__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_15__G2_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9373\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8941\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_571\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9492\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_0_14_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcccccccf0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_14__G2_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9509\,
datae => N_33607_1,
datad => N_29071_1,
datac => N_33222_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11810_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_6_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00300000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_1\,
dataf => N_32972,
datae => N_33543,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_603\,
datac => N_33734_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_12_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000c0000000000")
port map (
combout => N_32982,
dataf => N_32982_1,
datae => N_33179,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_1_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_1\,
datae => N_32978,
datad => N_32982,
datac => N_32722_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_8_TZ\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_1_2_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cc000c0000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_1_2\(13),
dataf => N_32844_2,
datae => N_33543,
datad => N_33368_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_2_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cf0f0f0fc0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_6_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_1_2\(13),
datae => N_28492_1,
datad => N_32909_1,
datac => N_34325_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_3_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c3000000000000")
port map (
combout => N_32973,
dataf => N_28492_1,
datae => N_32738_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_4_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_5\,
dataf => N_32976,
datae => N_32973,
datad => N_32970,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_16_0\(6),
datab => N_32956_I);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_3_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_8_0\,
dataf => N_32974,
datae => N_32844_3,
datad => N_32722_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_0_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff3000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_12\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_8_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_5\,
datad => N_32844_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_6_TZ\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_12\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_7\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_6_1\,
datac => N_34334,
datab => N_32981);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_0_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffcccf000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1079\,
datae => N_33794,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9503\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1607\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_811\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff0fc00cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8714\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1685\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9486\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_473\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9498\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1672\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8714\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_4\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_544\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_4_RNI79SG_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffc0ff00ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_0\,
dataf => N_32738_1,
datae => N_32844_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1049\,
datac => N_32762_I,
datab => N_33984_2);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_5_0_A2_RNI35C86_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000fc3c00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_4\,
dataf => N_32782_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_473\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9525\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_A2_25_RNI4EPKB_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff3f00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_15\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1044\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1768\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_7_RNI0FUUM_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_15\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_14\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8834\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_4\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_3_0_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c0000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_3_0\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_9_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cc0000000000000")
port map (
combout => N_33031,
dataf => N_34329_1,
datae => N_28652_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_4_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfc0000000000000")
port map (
combout => N_33026,
dataf => N_33297_1,
datae => N_32908_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff30000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_0\,
dataf => N_33026,
datae => N_28634_1,
datad => N_29262_1,
datac => N_33004,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_10\,
dataf => N_32848,
datae => N_33028,
datad => N_33024,
datac => N_33032,
datab => N_33023);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff8")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_10\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_8\,
datad => N_33021,
datac => N_33022,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_3_0\(4),
dataa => N_33010);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffc0c0c0ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2_1\,
dataf => N_34263_2,
datae => N_29071_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9490\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_1__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9349\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8631\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_0\(8),
datac => N_33794,
datab => N_28222_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_3_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00c000c000c00000")
port map (
combout => N_33780,
dataf => N_34254_1,
datae => N_32789_2,
datad => N_33111,
datac => N_32738_1_0,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_6_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000030000000")
port map (
combout => N_33783,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datae => N_32861_1,
datad => N_33140_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_1_RNIPA2E3_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00003000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_0\,
dataf => N_33778,
datae => N_29071_1,
datad => N_33140_1,
datac => N_34254_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_4_0_RNI93AB5_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffff030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_0\,
datae => N_33777,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A9_4_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffa080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_3\,
datad => N_33794,
datac => N_29262_1,
datab => N_33795,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_O2_11_RNI1VEE5_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff00ff000000ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_770\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_0_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0000000c000000")
port map (
combout => N_34039,
dataf => N_32861_1,
datae => N_32738_2,
datad => N_32738_1_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_3_RNIQ01Q2_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff30000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_4\,
dataf => N_34042,
datae => N_32723_1,
datad => N_33140_1,
datac => N_32818_I,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_6_1_RNIEPGN3_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff000000ff303030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_16_0\(6),
datad => N_34055_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_6_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_10_RNI56303_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00000030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_1\,
dataf => N_34049,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\,
datad => N_33140_1,
datac => N_28492_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O23_2_RNICMOL4_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00003000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
datad => N_32727_1,
datac => N_34024,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_0_RNIOC2PD1_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_17\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_16\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_6\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_5\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A32_6_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3cc3000000000000")
port map (
combout => N_33130,
dataf => N_29653_1,
datae => N_28211_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A32_3_1_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000c030f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A32_3_1\(57),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_604\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A32_2_0_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000f000f0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A32_2_0\(57),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_8_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0003000000000000")
port map (
combout => N_32978,
dataf => N_32844_3,
datae => N_28492_1,
datad => N_33368_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff003000f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_10\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1697\,
datae => N_29653_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_797\,
datac => N_32840_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A14_5_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c00000000000000")
port map (
combout => N_32843,
dataf => N_28634_1,
datae => N_29071_1,
datad => N_32722_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff30000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_1\,
dataf => N_32843,
datae => N_28634_1,
datad => N_33004,
datac => N_33146_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_1\,
datae => N_32844,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_797\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_3_1\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A14_4_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c300000000000000")
port map (
combout => N_32842,
dataf => N_32979_1,
datae => N_32738_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A14_9_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000003000000000")
port map (
combout => N_32847,
dataf => N_33140_1,
datae => N_33004,
datad => N_32818_I,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff000c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_3\,
dataf => N_32847,
datae => N_28857_1,
datad => N_32821,
datac => N_53933,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_10\,
datac => N_32848,
datab => N_32838);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_0_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000c0000")
port map (
combout => N_34255,
dataf => N_33368_1,
datae => N_32786_1,
datad => N_28261_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84));
\GRLFPC2_0_R_I_EXC_RNO_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000003000")
port map (
combout => \GRLFPC2_0.R.I.EXC_2_0_1__G2\,
dataf => \GRLFPC2_0.N_1438\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(40),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(38),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(41));
\GRLFPC2_0_R_I_EXC_RNO_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000cc00c000")
port map (
combout => \GRLFPC2_0.R.I.EXC_2_0_4__G2\,
dataf => \GRLFPC2_0.N_1438\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(40),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(38),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(41));
\GRLFPC2_0_R_A_RF2REN_RNO_0_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000fff")
port map (
combout => N_37405,
dataf => \GRLFPC2_0.N_951\,
datae => \GRLFPC2_0.RS1D_CNST\,
datad => \GRLFPC2_0.RS1V_0_SQMUXA\,
datac => N_78);
\GRLFPC2_0_R_A_RF2REN_RNO_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000f0003")
port map (
combout => N_37433,
dataf => \GRLFPC2_0.N_3477_1_I\,
datae => \GRLFPC2_0.N_2975\,
datad => N_37405,
datac => N_37362,
datab => \GRLFPC2_0.COMB.V.A.RF2REN_1_8055_I_A5_0_0\);
\GRLFPC2_0_R_A_RF1REN_RNO_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000003000f")
port map (
combout => N_37431,
dataf => \GRLFPC2_0.N_3477_1_I\,
datae => \GRLFPC2_0.N_2975\,
datad => N_37365_1,
datac => N_37362,
datab => \GRLFPC2_0.COMB.V.A.RF2REN_1_8055_I_A5_0_0\);
GRLFPC2_0_R_A_LD_RNO_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000c000000000")
port map (
combout => \GRLFPC2_0.R.A.LD_0_0_G1_3\,
dataf => \GRLFPC2_0.N_45\,
datae => N_75,
datad => N_74,
datac => N_84,
datab => N_83);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_D_108_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff000f0ffcc00cc")
port map (
combout => N_59001,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(108),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datac => \GRLFPC2_0.FPO.FRAC\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_D_109_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff000f0ffcc00cc")
port map (
combout => N_59000,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(109),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datac => \GRLFPC2_0.FPO.FRAC\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000003f003333ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2_16_TZ\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
GRLFPC2_0_R_X_FPOP_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
combout => \GRLFPC2_0.R.X.FPOP_0_0_G1\,
dataf => \GRLFPC2_0.R.M.FPOP\,
datae => N_294,
datad => N_295);
GRLFPC2_0_R_X_LD_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
combout => \GRLFPC2_0.R.X.LD_0_0_G1\,
dataf => \GRLFPC2_0.R.M.LD\,
datae => N_294,
datad => N_295);
GRLFPC2_0_R_M_AFSR_RET_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.R.M.AFSR_RET_0_0_G1\,
dataf => \GRLFPC2_0.N_1830_O\,
datae => \GRLFPC2_0.R.A.AFSR_O\);
GRLFPC2_0_R_M_AFQ_RET_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.R.M.AFQ_RET_0_0_G1\,
dataf => \GRLFPC2_0.N_1830_O\,
datae => \GRLFPC2_0.R.A.AFQ_O\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4459\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_53526,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(260));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_53503,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(261));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_53480,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(307));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_53457,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(308));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_53434,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(309));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_53416,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(310));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_21_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_53329,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(294));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_20_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_53306,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(295));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_53283,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(296));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_53260,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(297));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_53237,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(298));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_16_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_53214,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(299));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_15_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_53191,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(300));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_14_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_53168,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(301));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_53145,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(302));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_53122,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(303));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_53099,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(304));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_53076,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(305));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_9_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_53053,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(306));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_60_Z_1_SUM_0_0_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0f0ff00ff0f0f0")
port map (
combout => N_53048,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1274_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_53008,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(259));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_52985,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(279));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_35_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_52962,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(280));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_52939,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(281));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_52916,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(282));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_52893,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(283));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_52870,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(284));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_30_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_52847,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(285));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_52824,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(286));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_52801,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(287));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_52778,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(288));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_52755,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(289));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_52732,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(290));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_52709,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(291));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_23_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_52686,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(292));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_22_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_52663,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(293));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_52640,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(264));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_52617,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(265));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_52594,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(266));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_52571,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(267));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_52548,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(268));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_46_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_52525,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(269));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_45_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_52502,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(270));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_44_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_52479,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(271));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_43_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_52456,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(272));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_52433,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(273));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_41_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_52410,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(274));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_40_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_52387,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(275));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_52364,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(276));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff00ffffff00")
port map (
combout => N_52341,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(277));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_37_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_52318,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(278));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_52295,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(262));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_0_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => N_52272,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(263));
GRLFPC2_0_COMB_FPDECODE_RS1D5_0_A2_1_RNIGBRH: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3f3f00ff00000000")
port map (
combout => \GRLFPC2_0.COMB.V.A.RF2REN_1_8055_I_A5_0_0\,
dataf => \GRLFPC2_0.N_951\,
datae => N_72,
datad => \GRLFPC2_0.RS1D_CNST\,
datac => \GRLFPC2_0.COMB.FPDECODE.RS1D5_1\,
datab => \GRLFPC2_0.COMB.FPDECODE.RS1D5_0_A2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_233_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f3000000c000")
port map (
combout => N_37423,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(11),
datae => \GRLFPC2_0.FPI.LDOP_1_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7920_I_1_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIHKHD_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7920_I_1_1\,
dataf => \GRLFPC2_0.R.MK.RST2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datad => N_11);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_232_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000cf000000c000")
port map (
combout => N_37424,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(12),
datae => \GRLFPC2_0.FPI.LDOP_1_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7920_I_1_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(245));
GRLFPC2_0_COMB_V_STATE12: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c0ffffff00000000")
port map (
combout => \GRLFPC2_0.N_1015\,
dataf => \GRLFPC2_0.COMB.V.STATE12_0\,
datae => \GRLFPC2_0.COMB.UN1_MEXC_1\,
datad => \GRLFPC2_0.COMB.UN1_MEXC_0\,
datac => \GRLFPC2_0.R.FSR.TEM\(2),
datab => \GRLFPC2_0.R.I.EXC\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_5_S_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_A2_5_S\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1846\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_A2_14_S\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_492\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_2_3_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000003000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_A2_2_3\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1855\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1769\,
datad => N_32738_1_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83),
datab => N_59);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_2_3_RNIOL3L3_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000f03")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_TZ_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_A2_2_3\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_A2_5_S\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_4_TZ\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_A2_3_S\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_A2_14_S\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0f00000c000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_12\,
dataf => N_32982_1,
datae => N_33175,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f00000fff00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_4_TZ\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_6_1_0_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff0000ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_6_1_0\(51),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_7_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cfc0c0c0c0c0c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_8_TZ\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_5_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c030000ccc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_6_TZ\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3000300030303000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_13\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_719\,
datae => N_28261_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_32_1\(27),
datac => N_33984_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_3_RNISRAD4: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffccc0fcc0fccc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_317__G1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1281_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7035\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7034\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_316_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffccc0fcc0fccc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_316__G1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1281_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7035\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7051\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_CIN_3_RNI3QEC1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0c0fcc0fcf000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_318__G1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1281_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14_141_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_14\(141),
dataf => N_53995,
datae => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(143));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14_171_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_14\(171),
dataf => N_53995,
datae => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_O2_10_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff30ffffff3033")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_403\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1730\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1566\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856\,
datac => N_33652_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(66));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_O2_4_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffff0ff30")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1855\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_O2_4_0\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_743\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1540\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1839\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_429\);
GRLFPC2_0_FPCO_HOLDN_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => CPO_HOLDNZ,
dataf => \GRLFPC2_0.R.MK.HOLDN1\,
datae => \GRLFPC2_0.R.MK.HOLDN2\);
\GRLFPC2_0_COMB_DBGDATA_4_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff00f0f0")
port map (
combout => CPO_DBG_DATAZ(29),
dataf => N_400,
datae => N_401,
datad => N_695,
datac => N_631);
GRLFPC2_0_COMB_UN1_FPCI_4: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00ff0000")
port map (
combout => \GRLFPC2_0.COMB.UN1_FPCI_4\,
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS2\(0),
datad => \GRLFPC2_0.R.A.RS2D\);
\GRLFPC2_0_R_I_EXC_0_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000048c8c8c")
port map (
combout => \GRLFPC2_0.R.I.EXC_MB\(0),
dataf => \GRLFPC2_0.N_1438\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_28\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_27\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4664\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4662\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\);
\GRLFPC2_0_COMB_DBGDATA_4_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff00f0f0")
port map (
combout => CPO_DBG_DATAZ(12),
dataf => N_400,
datae => N_401,
datad => N_678,
datac => N_614);
\GRLFPC2_0_COMB_DBGDATA_4_15_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff00f0f0")
port map (
combout => CPO_DBG_DATAZ(15),
dataf => N_400,
datae => N_401,
datad => N_681,
datac => N_617);
GRLFPC2_0_R_A_AFQ_RET_2_RNIMUGP: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000f")
port map (
combout => \GRLFPC2_0.N_202\,
dataf => \GRLFPC2_0.FPCI_O\(0),
datae => \GRLFPC2_0.COMB.LOCKGEN.LOCKI_O\,
datad => \GRLFPC2_0.FPCI_O\(74),
datac => \GRLFPC2_0.FPCI_O\(73));
GRLFPC2_0_COMB_UN1_R_A_RS1_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000ff00")
port map (
combout => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
dataf => \GRLFPC2_0.N_1841\,
datae => \GRLFPC2_0.R.A.RS1D\,
datad => \GRLFPC2_0.R.A.RS1\(0));
GRLFPC2_0_COMB_V_E_STDATA2_0_O2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000ffff")
port map (
combout => \GRLFPC2_0.N_91\,
dataf => N_155,
datae => N_154);
GRLFPC2_0_COMB_UN1_R_A_RS1_1_0_O2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000ffff")
port map (
combout => \GRLFPC2_0.N_90\,
dataf => \GRLFPC2_0.R.STATE_O\(1),
datae => \GRLFPC2_0.R.STATE_O\(0));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_20_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000f0f0")
port map (
combout => \GRLFPC2_0.N_3103\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => N_686,
datac => N_622);
\GRLFPC2_0_COMB_DBGDATA_4_20_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff00f0f0")
port map (
combout => CPO_DBG_DATAZ(20),
dataf => N_400,
datae => N_401,
datad => N_686,
datac => N_622);
\GRLFPC2_0_COMB_DBGDATA_4_21_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff00f0f0")
port map (
combout => CPO_DBG_DATAZ(21),
dataf => N_400,
datae => N_401,
datad => N_687,
datac => N_623);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff00fffff0f0")
port map (
combout => \GRLFPC2_0.N_3101\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => N_684,
datac => N_620);
\GRLFPC2_0_COMB_DBGDATA_4_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffff00f0f0")
port map (
combout => CPO_DBG_DATAZ(17),
dataf => N_400,
datae => N_401,
datad => N_683,
datac => N_619);
\GRLFPC2_0_COMB_DBGDATA_4_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffff00f0f0")
port map (
combout => CPO_DBG_DATAZ(18),
dataf => N_400,
datae => N_401,
datad => N_684,
datac => N_620);
GRLFPC2_0_COMB_ANNULFPU_1_U_0_A3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000000000")
port map (
combout => \GRLFPC2_0.N_3491\,
dataf => \GRLFPC2_0.R.M.FPOP\,
datae => N_294,
datad => N_295);
GRLFPC2_0_WRADDR_1_SQMUXA: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f0ffffff")
port map (
combout => \GRLFPC2_0.WRADDR_1_SQMUXA\,
dataf => \GRLFPC2_0.N_1243\,
datae => \GRLFPC2_0.R.X.FPOP\,
datad => \GRLFPC2_0.R.I.V\,
datac => \GRLFPC2_0.R.I.EXEC\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_258_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cf3fffff30c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_258__N_5_I\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8_0\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6961\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_173_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0c000ccccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(173),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(173));
GRLFPC2_0_R_X_AFSR_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000f0000")
port map (
combout => \GRLFPC2_0.R.X.AFSR_0_0_G1\,
dataf => \GRLFPC2_0.N_1829_O\,
datae => \GRLFPC2_0.R.E.AFSR_O\,
datad => N_294,
datac => N_295);
GRLFPC2_0_R_X_AFQ_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000f0000")
port map (
combout => \GRLFPC2_0.R.X.AFQ_0_0_G1\,
dataf => \GRLFPC2_0.N_1829_O\,
datae => \GRLFPC2_0.R.E.AFQ_O\,
datad => N_294,
datac => N_295);
\GRLFPC2_0_R_I_CC_RNO_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff000000f000")
port map (
combout => \GRLFPC2_0.R.I.CC_0_0_0__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(40),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(13));
\GRLFPC2_0_R_I_CC_RNO_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff0000000f00")
port map (
combout => \GRLFPC2_0.R.I.CC_0_0_1__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(40),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(13));
GRLFPC2_0_R_I_PC_RET_60_RNI7KV4: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => N_13);
\GRLFPC2_0_R_FSR_FCC_RNO_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfc0cfc0cfcfc0c0")
port map (
combout => \GRLFPC2_0.R.FSR.FCC_0_0_1__G1\,
dataf => \GRLFPC2_0.N_1133\,
datae => \GRLFPC2_0.N_3227\,
datad => \GRLFPC2_0.R.I.CC\(1),
datac => \GRLFPC2_0.N_1517\,
datab => N_417);
\GRLFPC2_0_R_FSR_FCC_RNO_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfc0cfc0cfcfc0c0")
port map (
combout => \GRLFPC2_0.R.FSR.FCC_0_0_0__G1\,
dataf => \GRLFPC2_0.N_1133\,
datae => \GRLFPC2_0.N_3226\,
datad => \GRLFPC2_0.R.I.CC\(0),
datac => \GRLFPC2_0.N_1517\,
datab => N_416);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_45_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10089\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(45),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9969\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_45_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00ffff0f0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(45),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(45),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10207\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3c3f0c033033000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10018\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_3_I\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10103\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(31),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9983\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcc00ccf0f0f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9989\,
dataf => \GRLFPC2_0.FPI.LDOP_0_1\,
datae => \GRLFPC2_0.FPI.OP2\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(141),
datab => N_727);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cff0c00fcfffc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10109\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(25),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9989\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cff0c00fcfffc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10130\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10010\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10011\,
dataf => \GRLFPC2_0.FPI.LDOP_0_0\,
datae => \GRLFPC2_0.FPI.OP2\(54),
datad => \GRLFPC2_0.FPI.OP2\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(119));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cff0c00fcfffc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10131\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10011\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffccfcc33300300")
port map (
combout => N_54046,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(26),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00fff00f0fffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(25),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(25),
datae => N_54046,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff0ffff0ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(53),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(54),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"d9c8fbea51407362")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10019\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(55),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10035\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(39),
datae => \GRLFPC2_0.FPO.FRAC\(18),
datad => \GRLFPC2_0.FPO.FRAC\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_35_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10039\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(35),
datae => \GRLFPC2_0.FPO.FRAC\(22),
datad => \GRLFPC2_0.FPO.FRAC\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10040\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(34),
datae => \GRLFPC2_0.FPO.FRAC\(23),
datad => \GRLFPC2_0.FPO.FRAC\(22),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10045\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(29),
datae => \GRLFPC2_0.FPO.FRAC\(28),
datad => \GRLFPC2_0.FPO.FRAC\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10046\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(28),
datae => \GRLFPC2_0.FPO.FRAC\(29),
datad => \GRLFPC2_0.FPO.FRAC\(28),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbf8cbc83b380b08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10048\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(26),
datae => \GRLFPC2_0.FPO.FRAC\(30),
datad => \GRLFPC2_0.FPO.FRAC\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbf8cbc83b380b08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10049\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(25),
datae => \GRLFPC2_0.FPO.FRAC\(31),
datad => \GRLFPC2_0.FPO.FRAC\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_75_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0fff000ccffcc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(75),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.FPI.OP1\(37),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_674,
datab => N_610);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_72_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff000f0ffcc00cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(72),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.FPI.OP1\(43),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_674,
datab => N_610);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_69_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0fff000ccffcc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(69),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.FPI.OP1\(43),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_680,
datab => N_616);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_66_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff000f0ffcc00cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(66),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.FPI.OP1\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_680,
datab => N_616);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_63_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0fff000ccffcc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(63),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.FPI.OP1\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_686,
datab => N_622);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_254_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfffcf00c0ffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10520\,
dataf => \GRLFPC2_0.FPO.EXP\(4),
datae => \GRLFPC2_0.FPO.EXP\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(241));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_64_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff000f0ffcc00cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(64),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.FPI.OP1\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_682,
datab => N_618);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_255_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfffcf00c0ffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10519\,
dataf => \GRLFPC2_0.FPO.EXP\(3),
datae => \GRLFPC2_0.FPO.EXP\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0d0c0c0c0d0c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10934\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7786\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM12\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10931\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"faffccfffa00cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10934\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10007\,
dataf => \GRLFPC2_0.FPI.LDOP_0_1\,
datae => \GRLFPC2_0.FPI.OP2\(50),
datad => \GRLFPC2_0.FPI.OP2\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(123));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cff0c00fcfffc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10127\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10007\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_20_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbf8cbc83b380b08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10054\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(20),
datae => \GRLFPC2_0.FPO.FRAC\(36),
datad => \GRLFPC2_0.FPO.FRAC\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_4_0_RNIPHTL2_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33f0cc00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7034\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6961\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_258_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00fff00ff00fff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8_0\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1281_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7035\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_4_0_RNI8FMJ1_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fccf000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7051\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6961\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bcb0bf838c808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10074\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_175__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbf8cbc83b380b08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10047\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(27),
datae => \GRLFPC2_0.FPO.FRAC\(29),
datad => \GRLFPC2_0.FPO.FRAC\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10032\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(42),
datae => \GRLFPC2_0.FPO.FRAC\(15),
datad => \GRLFPC2_0.FPO.FRAC\(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_43_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10031\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(43),
datae => \GRLFPC2_0.FPO.FRAC\(14),
datad => \GRLFPC2_0.FPO.FRAC\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_41_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10033\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(41),
datae => \GRLFPC2_0.FPO.FRAC\(16),
datad => \GRLFPC2_0.FPO.FRAC\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10108\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(26),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9988\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcf3f00f0c0300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(26),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(28),
datae => N_53989,
datad => N_53977,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcff3000fc0030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(2),
datae => N_53982,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datac => N_53942,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10027\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(47),
datae => \GRLFPC2_0.FPO.FRAC\(10),
datad => \GRLFPC2_0.FPO.FRAC\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_44_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10030\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(44),
datae => \GRLFPC2_0.FPO.FRAC\(13),
datad => \GRLFPC2_0.FPO.FRAC\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10084\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(50),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9964\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10096\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(38),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9976\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(50),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_14_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10000\,
dataf => \GRLFPC2_0.FPI.LDOP_0_1\,
datae => \GRLFPC2_0.FPI.OP2\(43),
datad => \GRLFPC2_0.FPI.OP2\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(130));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_14_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30ff3000fcfffc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10120\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(14),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10000\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_14_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(14),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(43),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(15),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10107\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(27),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9987\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => N_54039,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(27),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(30),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(28),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00fff00f0fffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(27),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(27),
datae => N_54039,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_44_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10090\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(44),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9970\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_44_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f33fff00c00ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(44),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(13),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_45_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10029\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(45),
datae => \GRLFPC2_0.FPO.FRAC\(12),
datad => \GRLFPC2_0.FPO.FRAC\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffccfff000cc00f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(28),
dataf => N_53963,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffccfcc33300300")
port map (
combout => N_54042,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(29),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(30),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(28),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00fff00f0fffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(28),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(28),
datae => N_54042,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10106\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(28),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9986\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbf8cbc83b380b08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10055\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(19),
datae => \GRLFPC2_0.FPO.FRAC\(37),
datad => \GRLFPC2_0.FPO.FRAC\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10003\,
dataf => \GRLFPC2_0.FPI.LDOP_0_1\,
datae => \GRLFPC2_0.FPI.OP2\(46),
datad => \GRLFPC2_0.FPI.OP2\(43),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(127));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cff0c00fcfffc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10123\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(11),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10003\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f33fff00c00ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(11),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(46),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10087\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(47),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9967\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ff333cc0cc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(10),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(10),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(47),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10004\,
dataf => \GRLFPC2_0.FPI.LDOP_0_1\,
datae => \GRLFPC2_0.FPI.OP2\(47),
datad => \GRLFPC2_0.FPI.OP2\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(126));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cff0c00fcfffc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10124\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(10),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10004\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00cfc03f30fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9783\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10197\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_248_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10512\,
dataf => \GRLFPC2_0.FPO.EXP\(10),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_246_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10514\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(12),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_256_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfffcf00c0ffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10518\,
dataf => \GRLFPC2_0.FPO.EXP\(2),
datae => \GRLFPC2_0.FPO.EXP\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_253_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfffcf00c0ffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10521\,
dataf => \GRLFPC2_0.FPO.EXP\(5),
datae => \GRLFPC2_0.FPO.EXP\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(240));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_250_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfffcf00c0ffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10524\,
dataf => \GRLFPC2_0.FPO.EXP\(8),
datae => \GRLFPC2_0.FPO.EXP\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(237));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_CIN_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33f0cc00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6961\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fccf000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6583\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_CIN_3_RNI3QEC1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f00f3cc33cc30ff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1281_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bf838cb0bc808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10072\,
dataf => \GRLFPC2_0.FPO.FRAC\(54),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_176__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00fff0ff0fffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(52),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f33fff00c00ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(52),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10009\,
dataf => \GRLFPC2_0.FPI.LDOP_0_0\,
datae => \GRLFPC2_0.FPI.OP2\(52),
datad => \GRLFPC2_0.FPI.OP2\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(121));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cff0c00fcfffc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10129\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10009\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10100\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9980\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0cc00ccffcc0fcc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9805\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(24),
datae => N_54033,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(34),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(23),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(35),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcffccc33033000")
port map (
combout => N_54033,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10025\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(49),
datae => \GRLFPC2_0.FPO.FRAC\(8),
datad => \GRLFPC2_0.FPO.FRAC\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ccf0cc0fccffcc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9789\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10203\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3fcf0ff030c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(49),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(49),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_45_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cc0cc000ff3ff333")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10207\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(45),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(46),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00cfc03f30fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9781\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10195\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(115),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfc00f00fff03f30")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9782\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(1),
datae => N_54031,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN5_SHDVAR: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffcfcff33fc30")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN5_SHDVAR\,
dataf => N_53909,
datae => N_53915,
datad => N_53913,
datac => N_53916,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN38_SHDVAR_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN38_SHDVAR_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN20_SHDVAR: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccccccccccccc0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN20_SHDVAR\,
dataf => N_53916,
datae => N_53915,
datad => N_53917,
datac => N_53914,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_2_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000003000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(57),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN5_SHDVAR\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN20_SHDVAR\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN40_SHDVAR\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10023\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(51),
datae => \GRLFPC2_0.FPO.FRAC\(6),
datad => \GRLFPC2_0.FPO.FRAC\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f33fff00c00ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(38),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(19),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10010\,
dataf => \GRLFPC2_0.FPI.LDOP_0_0\,
datae => \GRLFPC2_0.FPI.OP2\(53),
datad => \GRLFPC2_0.FPI.OP2\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(120));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcf3f00f0c0300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(7),
datae => N_53948,
datad => N_53935,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffccfcc33300300")
port map (
combout => N_54028,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcf3f00f0c0300")
port map (
combout => N_53994,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00fff00f0fffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(7),
dataf => N_53994,
datae => N_54028,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_30_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10044\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(30),
datae => \GRLFPC2_0.FPO.FRAC\(27),
datad => \GRLFPC2_0.FPO.FRAC\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3fcf00f030c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(11),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(13),
datae => N_53955,
datad => N_53974,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff033f0ccf000f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(34),
dataf => N_53964,
datae => N_53961,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10105\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(29),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9985\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f33fff00c00ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(31),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(26),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3fcf0ff030c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(29),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(29),
datae => N_53957,
datad => N_53966,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_40_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10094\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(40),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9974\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_40_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(40),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(41),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_40_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10034\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(40),
datae => \GRLFPC2_0.FPO.FRAC\(17),
datad => \GRLFPC2_0.FPO.FRAC\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_43_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10091\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(43),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9971\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_43_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f33fff00c00ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(43),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(14),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(43),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_45_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3fff0cff3f000c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(45),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(45),
datae => N_53972,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10021\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(53),
datae => \GRLFPC2_0.FPO.FRAC\(4),
datad => \GRLFPC2_0.FPO.FRAC\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10022\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(52),
datae => \GRLFPC2_0.FPO.FRAC\(5),
datad => \GRLFPC2_0.FPO.FRAC\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10080\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(54),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9960\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10024\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(50),
datae => \GRLFPC2_0.FPO.FRAC\(7),
datad => \GRLFPC2_0.FPO.FRAC\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10026\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(48),
datae => \GRLFPC2_0.FPO.FRAC\(9),
datad => \GRLFPC2_0.FPO.FRAC\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_46_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10028\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(46),
datae => \GRLFPC2_0.FPO.FRAC\(11),
datad => \GRLFPC2_0.FPO.FRAC\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10086\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(48),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9966\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ccf033f000f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(50),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcffccc33033000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10203\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(50),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ff333cc0cc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10204\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(48),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3fcf00f030c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(48),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(47),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcffccc33033000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(48),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(48),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00ffff0f0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(48),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(48),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10204\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10020\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(54),
datae => \GRLFPC2_0.FPO.FRAC\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIKTCN2_315_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f0ffffffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1_1\,
dataf => N_53999,
datae => N_53997,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(315));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN36_STKGEN_0_0_RNI3CM9J: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"eddfefdefdfffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN25_NOTPROP\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN36_STKGEN_0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SCLSBS_2\(0),
datac => N_54002,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5458\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f00ff000000f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10017\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f33fff00c00ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(36),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(21),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10098\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(36),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9978\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10095\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(39),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9975\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_40_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf3f0ff0c03000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(40),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(40),
datae => N_53986,
datad => N_53988,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff033f0ccf000f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(39),
dataf => N_53970,
datae => N_53971,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(39),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(39),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(18),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(40),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53916,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffccfcc33300300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(57),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(55),
datae => N_53913,
datad => N_53916,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(8),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10066\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(8),
datae => \GRLFPC2_0.FPO.FRAC\(49),
datad => \GRLFPC2_0.FPO.FRAC\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbf8cbc83b380b08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10067\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(7),
datae => \GRLFPC2_0.FPO.FRAC\(49),
datad => \GRLFPC2_0.FPO.FRAC\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bcb0bf838c808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10069\,
dataf => \GRLFPC2_0.FPO.FRAC\(52),
datae => \GRLFPC2_0.FPO.FRAC\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bf838cb0bc808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10070\,
dataf => \GRLFPC2_0.FPO.FRAC\(52),
datae => \GRLFPC2_0.FPO.FRAC\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ffcc00f000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(7),
dataf => N_53955,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf3f0ff0c03000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(6),
datae => N_53981,
datad => N_53980,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => N_54021,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10008\,
dataf => \GRLFPC2_0.FPI.LDOP_0_1\,
datae => \GRLFPC2_0.FPI.OP2\(51),
datad => \GRLFPC2_0.FPI.OP2\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(122));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30ff3000fcfffc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10128\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10008\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_21_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbf8cbc83b380b08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10053\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(21),
datae => \GRLFPC2_0.FPO.FRAC\(35),
datad => \GRLFPC2_0.FPO.FRAC\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0cfc03f300f00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(3),
dataf => N_53948,
datae => N_53935,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f33fff00c00ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(55),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_80_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0fff000ccffcc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(80),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.FPI.OP1\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_669,
datab => N_605);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_77_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff000f0ffcc00cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(77),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.FPI.OP1\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_669,
datab => N_605);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_65_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0fff000ccffcc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(65),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.FPI.OP1\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_684,
datab => N_620);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff000f0ffcc00cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(62),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.FPI.OP1\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_684,
datab => N_620);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_14_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf3f0ff0c03000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(14),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(14),
datae => N_53946,
datad => N_53947,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcffccc33033000")
port map (
combout => N_54022,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(14),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33c30cfc30c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(13),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(11),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(12),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00fff00f0fffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(13),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(13),
datae => N_54022,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10001\,
dataf => \GRLFPC2_0.FPI.LDOP_0_1\,
datae => \GRLFPC2_0.FPI.OP2\(44),
datad => \GRLFPC2_0.FPI.OP2\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(129));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30ff3000fcfffc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10121\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(13),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10001\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbf8cbc83b380b08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10064\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(10),
datae => \GRLFPC2_0.FPO.FRAC\(46),
datad => \GRLFPC2_0.FPO.FRAC\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_37_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10097\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(37),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9977\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_22_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9992\,
dataf => \GRLFPC2_0.FPI.LDOP_0_1\,
datae => \GRLFPC2_0.FPI.OP2\(35),
datad => \GRLFPC2_0.FPI.OP2\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(138));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_22_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30ff3000fcfffc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10112\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(22),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9992\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0ff000cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9995\,
dataf => \GRLFPC2_0.FPI.LDOP_0_1\,
datae => \GRLFPC2_0.FPI.OP2\(35),
datad => \GRLFPC2_0.FPI.OP2\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(135));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"30ff3000fcfffc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10115\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(19),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9995\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_15_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9999\,
dataf => \GRLFPC2_0.FPI.LDOP_0_1\,
datae => \GRLFPC2_0.FPI.OP2\(42),
datad => \GRLFPC2_0.FPI.OP2\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(131));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_15_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cff0c00fcfffc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10119\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(15),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9999\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10002\,
dataf => \GRLFPC2_0.FPI.LDOP_0_1\,
datae => \GRLFPC2_0.FPI.OP2\(45),
datad => \GRLFPC2_0.FPI.OP2\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(128));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cff0c00fcfffc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10122\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(12),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10002\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_9_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10005\,
dataf => \GRLFPC2_0.FPI.LDOP_0_1\,
datae => \GRLFPC2_0.FPI.OP2\(48),
datad => \GRLFPC2_0.FPI.OP2\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(125));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_9_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cff0c00fcfffc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10125\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(9),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10005\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_37_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00fcfcff003030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(37),
dataf => N_53970,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(39),
datac => N_53962,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_37_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(37),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(20),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffccfcc33300300")
port map (
combout => N_54017,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(20),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(21),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00fff00f0fffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(19),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(19),
datae => N_54017,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_15_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf3f0ff0c03000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(15),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(15),
datae => N_53979,
datad => N_53978,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_15_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f33fff00c00ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(15),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(42),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(15),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffccfff000cc00f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(13),
dataf => N_53978,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcf3f00f0c0300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(12),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(14),
datae => N_53947,
datad => N_53981,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ff333cc0cc000")
port map (
combout => N_54015,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(12),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3cfc33c300c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(12),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(11),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(10),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00fff00f0fffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(12),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(12),
datae => N_54015,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf3f0ff0c03000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(10),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(10),
datae => N_53947,
datad => N_53981,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcc00ccf0f0f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9990\,
dataf => \GRLFPC2_0.FPI.LDOP_0_1\,
datae => \GRLFPC2_0.FPI.OP2\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(140),
datab => N_728);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cff0c00fcfffc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10110\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(24),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9990\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ffcc00f000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(27),
dataf => N_53957,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => N_54013,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(24),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00fff00f0fffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(24),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(24),
datae => N_54013,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10102\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9982\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_30_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10104\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(30),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9984\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0fff0ccf033f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(32),
dataf => N_53964,
datae => N_53963,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ff333cc0cc000")
port map (
combout => N_54012,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53976,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53957,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3ffc000f300c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(31),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(33),
datae => N_53957,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datac => N_53966,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53963,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_30_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf3f0ff0c03000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(30),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(30),
datae => N_53964,
datad => N_53963,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_30_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f33fff00c00ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(30),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(27),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(30),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10092\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(42),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9972\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(42),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(15),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(43),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_41_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10093\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(41),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9973\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_35_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10099\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(35),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9979\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53952,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcf3f00f0c0300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(42),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(44),
datae => N_53986,
datad => N_53988,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53971,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_41_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3fcf00f030c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(41),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(43),
datae => N_53970,
datad => N_53971,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_41_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(41),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(16),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_15_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53988,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53961,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_21_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53964,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3fcf00f030c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(36),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(38),
datae => N_53964,
datad => N_53961,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_16_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53970,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_20_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53962,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_22_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53966,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_35_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcff30fffc003000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(35),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(35),
datae => N_53970,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datac => N_53962,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_35_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(35),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(22),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10081\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(53),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9961\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0cff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10082\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(52),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9962\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ff333cc0cc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ff333cc0cc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(52),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_46_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10088\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(46),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9968\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53973,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53972,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffc0fff300c000f3")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(49),
datae => N_53972,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_9_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53953,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53986,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_46_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcffccc33033000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10206\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(47),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(46),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_46_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00ffff0f0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(46),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(46),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10206\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_16_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcf3f00f0c0300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(16),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(18),
datae => N_53946,
datad => N_53947,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_16_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0000ff0000")
port map (
combout => N_54041,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(16),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_16_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfc00f00fff03f30")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9822\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(41),
datae => N_54041,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fcff30fffc003000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(51),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(51),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffccfcc33300300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(51),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(49),
datae => N_53888,
datad => N_53912,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf3f0ff0c03000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(51),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(51),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcf3f00f0c0300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(50),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(49),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ff333cc0cc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(51),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_I\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3030ff00fcfcff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(51),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9963\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_45_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33c30cfc30c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(45),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(43),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53915,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffccfcc33300300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(56),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(54),
datae => N_53909,
datad => N_53915,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53914,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0ff00ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8_I\(57),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10042\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(32),
datae => \GRLFPC2_0.FPO.FRAC\(25),
datad => \GRLFPC2_0.FPO.FRAC\(24),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_23_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbf8cbc83b380b08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10051\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(23),
datae => \GRLFPC2_0.FPO.FRAC\(33),
datad => \GRLFPC2_0.FPO.FRAC\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_22_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbf8cbc83b380b08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10052\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(22),
datae => \GRLFPC2_0.FPO.FRAC\(34),
datad => \GRLFPC2_0.FPO.FRAC\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbf8cbc83b380b08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10050\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(24),
datae => \GRLFPC2_0.FPO.FRAC\(32),
datad => \GRLFPC2_0.FPO.FRAC\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbf8cbc83b380b08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10061\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(13),
datae => \GRLFPC2_0.FPO.FRAC\(43),
datad => \GRLFPC2_0.FPO.FRAC\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_37_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcffccc33033000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(37),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(35),
datae => N_53892,
datad => N_53904,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_37_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3fcf0ff030c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(37),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(37),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fb3bcb0bf838c808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10071\,
dataf => \GRLFPC2_0.FPO.FRAC\(54),
datae => \GRLFPC2_0.FPO.FRAC\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10041\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(33),
datae => \GRLFPC2_0.FPO.FRAC\(24),
datad => \GRLFPC2_0.FPO.FRAC\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10043\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(31),
datae => \GRLFPC2_0.FPO.FRAC\(26),
datad => \GRLFPC2_0.FPO.FRAC\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10036\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(38),
datae => \GRLFPC2_0.FPO.FRAC\(19),
datad => \GRLFPC2_0.FPO.FRAC\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cff0c00fcfffc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10126\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10006\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53974,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_46_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53955,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_9_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccfff0ffcc00f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(9),
dataf => N_53948,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_9_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3fcf0ff030c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(9),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(9),
datae => N_53955,
datad => N_53974,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_45_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53981,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcf3f00f0c0300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(8),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(10),
datae => N_53981,
datad => N_53980,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(8),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(49),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53948,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9997\,
dataf => \GRLFPC2_0.FPI.LDOP_0_1\,
datae => \GRLFPC2_0.FPI.OP2\(40),
datad => \GRLFPC2_0.FPI.OP2\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(133));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cff0c00fcfffc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10117\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9997\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_40_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53978,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcf3f00f0c0300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(17),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(19),
datae => N_53979,
datad => N_53978,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33f33fff00c00ccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(17),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(40),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf3c0cf3c33000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(19),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(19),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfc00f00fff03f30")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9820\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(39),
datae => N_54005,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53956,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => N_54005,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(18),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(21),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53959,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccfff0ffcc00f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(18),
dataf => N_53959,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3fcf0ff030c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(18),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(18),
datae => N_53946,
datad => N_53945,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3cfc33c300c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(24),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(23),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(22),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(24),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_23_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcc00ccf0f0f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9991\,
dataf => \GRLFPC2_0.FPI.LDOP_0_1\,
datae => \GRLFPC2_0.FPI.OP2\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(139),
datab => N_729);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_23_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cff0c00fcfffc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10111\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(23),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9991\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53989,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf3f0ff0c03000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(24),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(24),
datae => N_53989,
datad => N_53977,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53969,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_23_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(23),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(24),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_30_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3fcf00f030c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(30),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(29),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(30),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(28),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(28),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(28),
datae => N_53908,
datad => N_53890,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ccf0cf330c300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(28),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(28),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(26),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcff3c33c0c3000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(27),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(26),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffccfcc33300300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(26),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(24),
datae => N_53908,
datad => N_53890,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3cf330cf0cc300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(26),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(24),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(26),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33c30cfc30c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(25),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(23),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(24),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_37_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10037\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(37),
datae => \GRLFPC2_0.FPO.FRAC\(20),
datad => \GRLFPC2_0.FPO.FRAC\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_41_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53947,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_43_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(43),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(43),
datae => N_53892,
datad => N_53891,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ff333cc0cc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(42),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(42),
datae => N_53886,
datad => N_53885,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53917,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53909,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53912,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53911,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53913,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(53),
datae => N_53888,
datad => N_53912,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(47),
datae => N_53891,
datad => N_53882,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_46_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(46),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(46),
datae => N_53886,
datad => N_53922,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53922,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_44_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffccfcc33300300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(44),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(42),
datae => N_53886,
datad => N_53922,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_14_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53901,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_45_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffccfcc33300300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(45),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(43),
datae => N_53891,
datad => N_53882,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_46_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33c30cfc30c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(46),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(44),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(45),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10006\,
dataf => \GRLFPC2_0.FPI.LDOP_0_1\,
datae => \GRLFPC2_0.FPI.OP2\(49),
datad => \GRLFPC2_0.FPI.OP2\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(124));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3fcf00f030c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(36),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(35),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_35_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf3f0ff0c03000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(35),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(35),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53888,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_122_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_116_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23));
\GRLFPC2_0_RS1_1_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => RFI2_RD1ADDRZ(3),
dataf => \GRLFPC2_0.COMB.RS1_1\(4),
datae => N_405,
datad => N_398);
\GRLFPC2_0_COMB_V_E_STDATA_1_0_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcc3300fcfc3030")
port map (
combout => \GRLFPC2_0.N_3078\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.INST\(28),
datad => \GRLFPC2_0.FPCI_O\(311),
datac => \GRLFPC2_0.R.I.PC_O\(28),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_COMB_DBGDATA_4_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(10),
dataf => CPO_CCZ(0),
datae => N_400,
datad => N_401,
datac => N_676,
datab => N_612);
\GRLFPC2_0_COMB_DBGDATA_4_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(24),
dataf => \GRLFPC2_0.R.FSR.TEM\(1),
datae => N_400,
datad => N_401,
datac => N_690,
datab => N_626);
\GRLFPC2_0_COMB_DBGDATA_4_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(27),
dataf => \GRLFPC2_0.R.FSR.TEM\(4),
datae => N_400,
datad => N_401,
datac => N_693,
datab => N_629);
\GRLFPC2_0_COMB_WRDATA_4_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(10),
dataf => \GRLFPC2_0.R.I.RES\(39),
datae => \GRLFPC2_0.R.I.RES\(10),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(10),
dataf => N_416,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_376,
datab => \GRLFPC2_0.COMB.WRDATA_4\(10));
\GRLFPC2_0_COMB_WRDATA_4_23_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(23),
dataf => \GRLFPC2_0.R.I.RES\(52),
datae => \GRLFPC2_0.R.I.RES\(23),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_23_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(23),
dataf => N_429,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_389,
datab => \GRLFPC2_0.COMB.WRDATA_4\(23));
\GRLFPC2_0_COMB_WRDATA_4_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(55),
dataf => \GRLFPC2_0.R.I.RES\(52),
datae => \GRLFPC2_0.R.I.RES\(55),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(23),
dataf => N_429,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_389,
datab => \GRLFPC2_0.COMB.WRDATA_4\(55));
\GRLFPC2_0_COMB_DBGDATA_4_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(0),
dataf => \GRLFPC2_0.R.FSR.CEXC\(0),
datae => N_400,
datad => N_401,
datac => N_666,
datab => N_602);
\GRLFPC2_0_COMB_DBGDATA_4_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(3),
dataf => \GRLFPC2_0.R.FSR.CEXC\(3),
datae => N_400,
datad => N_401,
datac => N_669,
datab => N_605);
\GRLFPC2_0_COMB_DBGDATA_4_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(4),
dataf => \GRLFPC2_0.R.FSR.CEXC\(4),
datae => N_400,
datad => N_401,
datac => N_670,
datab => N_606);
\GRLFPC2_0_COMB_WRDATA_4_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(8),
dataf => \GRLFPC2_0.R.I.RES\(37),
datae => \GRLFPC2_0.R.I.RES\(8),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(8),
dataf => N_414,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_374,
datab => \GRLFPC2_0.COMB.WRDATA_4\(8));
\GRLFPC2_0_COMB_WRDATA_4_15_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(15),
dataf => \GRLFPC2_0.R.I.RES\(44),
datae => \GRLFPC2_0.R.I.RES\(15),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_15_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(15),
dataf => N_421,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_381,
datab => \GRLFPC2_0.COMB.WRDATA_4\(15));
\GRLFPC2_0_COMB_WRDATA_4_21_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(21),
dataf => \GRLFPC2_0.R.I.RES\(50),
datae => \GRLFPC2_0.R.I.RES\(21),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_21_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(21),
dataf => N_427,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_387,
datab => \GRLFPC2_0.COMB.WRDATA_4\(21));
\GRLFPC2_0_COMB_WRDATA_4_40_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(40),
dataf => \GRLFPC2_0.R.I.RES\(37),
datae => \GRLFPC2_0.R.I.RES\(40),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_40_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(8),
dataf => N_414,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_374,
datab => \GRLFPC2_0.COMB.WRDATA_4\(40));
\GRLFPC2_0_COMB_WRDATA_4_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(47),
dataf => \GRLFPC2_0.R.I.RES\(44),
datae => \GRLFPC2_0.R.I.RES\(47),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(15),
dataf => N_421,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_381,
datab => \GRLFPC2_0.COMB.WRDATA_4\(47));
\GRLFPC2_0_COMB_WRDATA_4_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(53),
dataf => \GRLFPC2_0.R.I.RES\(50),
datae => \GRLFPC2_0.R.I.RES\(53),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(21),
dataf => N_427,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_387,
datab => \GRLFPC2_0.COMB.WRDATA_4\(53));
\GRLFPC2_0_RS1_1_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => RFI2_RD1ADDRZ(1),
dataf => \GRLFPC2_0.COMB.RS1_1\(2),
datae => N_403,
datad => N_398);
\GRLFPC2_0_RS1_1_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => RFI2_RD1ADDRZ(2),
dataf => \GRLFPC2_0.COMB.RS1_1\(3),
datae => N_404,
datad => N_398);
\GRLFPC2_0_RS2_1_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => RFI2_RD2ADDRZ(0),
dataf => \GRLFPC2_0.COMB.RS2_1\(1),
datae => N_402,
datad => N_398);
\GRLFPC2_0_RS2_1_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => RFI2_RD2ADDRZ(1),
dataf => \GRLFPC2_0.COMB.RS2_1\(2),
datae => N_403,
datad => N_398);
\GRLFPC2_0_COMB_RS2_1_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000fffff0000000")
port map (
combout => \GRLFPC2_0.COMB.RS2_1\(3),
dataf => \GRLFPC2_0.R.A.RS2\(3),
datae => N_13,
datad => \GRLFPC2_0.N_951\,
datac => N_56);
\GRLFPC2_0_RS2_1_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => RFI2_RD2ADDRZ(2),
dataf => \GRLFPC2_0.COMB.RS2_1\(3),
datae => N_404,
datad => N_398);
\GRLFPC2_0_COMB_RS2_1_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000fffff0000000")
port map (
combout => \GRLFPC2_0.COMB.RS2_1\(4),
dataf => \GRLFPC2_0.R.A.RS2\(4),
datae => N_13,
datad => \GRLFPC2_0.N_951\,
datac => N_57);
\GRLFPC2_0_RS2_1_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => RFI2_RD2ADDRZ(3),
dataf => \GRLFPC2_0.COMB.RS2_1\(4),
datae => N_405,
datad => N_398);
\GRLFPC2_0_COMB_RF2REN_1_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0ccfffff0cc")
port map (
combout => RFI2_REN1Z,
dataf => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT\,
datae => N_398,
datad => N_13,
datac => \GRLFPC2_0.COMB.V.A.RF2REN_1\(1),
datab => \GRLFPC2_0.R.A.RF2REN\(1));
\GRLFPC2_0_COMB_RF1REN_1_0_0_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3f0ffff33003300")
port map (
combout => \GRLFPC2_0.N_3150\,
dataf => \GRLFPC2_0.N_3475\,
datae => \GRLFPC2_0.COMB.RS2_1\(0),
datad => \GRLFPC2_0.R.A.RF1REN\(2),
datac => \GRLFPC2_0.N_77_1\,
datab => N_13);
GRLFPC2_0_COMB_UN31_DEBUG_UNIT: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT\,
dataf => N_400,
datae => N_399);
\GRLFPC2_0_COMB_RF1REN_1_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0ccfffff0cc")
port map (
combout => RFI1_REN1Z,
dataf => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT\,
datae => N_398,
datad => N_13,
datac => \GRLFPC2_0.COMB.V.A.RF1REN_1\(1),
datab => \GRLFPC2_0.R.A.RF1REN\(1));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00fc30fc30")
port map (
combout => \GRLFPC2_0.N_3056\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.FPCI_O\(289),
datad => \GRLFPC2_0.R.I.INST\(6),
datac => \GRLFPC2_0.R.I.PC_O\(6),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_COMB_V_I_PC_1_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.R.I.PC\(7),
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.FPCI_O\(290),
datad => \GRLFPC2_0.R.I.PC_O\(7));
\GRLFPC2_0_COMB_DBGDATA_4_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(5),
dataf => \GRLFPC2_0.R.FSR.AEXC\(0),
datae => N_400,
datad => N_401,
datac => N_671,
datab => N_607);
\GRLFPC2_0_COMB_WRDATA_4_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(27),
dataf => \GRLFPC2_0.R.I.RES\(56),
datae => \GRLFPC2_0.R.I.RES\(27),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(27),
dataf => N_433,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_393,
datab => \GRLFPC2_0.COMB.WRDATA_4\(27));
\GRLFPC2_0_COMB_WRDATA_4_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(31),
dataf => \GRLFPC2_0.R.I.RES\(63),
datae => \GRLFPC2_0.R.I.RES\(31),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(31),
dataf => N_437,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_397,
datab => \GRLFPC2_0.COMB.WRDATA_4\(31));
\GRLFPC2_0_COMB_WRDATA_4_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(54),
dataf => \GRLFPC2_0.R.I.RES\(51),
datae => \GRLFPC2_0.R.I.RES\(54),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(22),
dataf => N_428,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_388,
datab => \GRLFPC2_0.COMB.WRDATA_4\(54));
\GRLFPC2_0_COMB_WRDATA_4_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(59),
dataf => \GRLFPC2_0.R.I.RES\(56),
datae => \GRLFPC2_0.R.I.RES\(59),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(27),
dataf => N_433,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_393,
datab => \GRLFPC2_0.COMB.WRDATA_4\(59));
\GRLFPC2_0_WRDATA_63_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(31),
dataf => N_437,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_397,
datab => \GRLFPC2_0.R.I.RES\(63));
\GRLFPC2_0_COMB_DBGDATA_4_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(8),
dataf => \GRLFPC2_0.R.FSR.AEXC\(3),
datae => N_400,
datad => N_401,
datac => N_674,
datab => N_610);
\GRLFPC2_0_COMB_DBGDATA_4_9_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(9),
dataf => \GRLFPC2_0.R.FSR.AEXC\(4),
datae => N_400,
datad => N_401,
datac => N_675,
datab => N_611);
\GRLFPC2_0_COMB_DBGDATA_4_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(11),
dataf => CPO_CCZ(1),
datae => N_400,
datad => N_401,
datac => N_677,
datab => N_613);
\GRLFPC2_0_COMB_WRDATA_4_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(62),
dataf => \GRLFPC2_0.R.I.RES\(59),
datae => \GRLFPC2_0.R.I.RES\(62),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(30),
dataf => N_436,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_396,
datab => \GRLFPC2_0.COMB.WRDATA_4\(62));
\GRLFPC2_0_COMB_DBGDATA_4_22_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(22),
dataf => \GRLFPC2_0.R.FSR.NONSTD\,
datae => N_400,
datad => N_401,
datac => N_688,
datab => N_624);
\GRLFPC2_0_COMB_WRDATA_4_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(0),
dataf => \GRLFPC2_0.R.I.RES\(29),
datae => \GRLFPC2_0.R.I.RES\(0),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(0),
dataf => N_406,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_366,
datab => \GRLFPC2_0.COMB.WRDATA_4\(0));
\GRLFPC2_0_COMB_WRDATA_4_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(2),
dataf => \GRLFPC2_0.R.I.RES\(31),
datae => \GRLFPC2_0.R.I.RES\(2),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(2),
dataf => N_408,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_368,
datab => \GRLFPC2_0.COMB.WRDATA_4\(2));
\GRLFPC2_0_COMB_WRDATA_4_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(3),
dataf => \GRLFPC2_0.R.I.RES\(32),
datae => \GRLFPC2_0.R.I.RES\(3),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(3),
dataf => N_409,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_369,
datab => \GRLFPC2_0.COMB.WRDATA_4\(3));
\GRLFPC2_0_COMB_WRDATA_4_22_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(22),
dataf => \GRLFPC2_0.R.I.RES\(51),
datae => \GRLFPC2_0.R.I.RES\(22),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_22_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(22),
dataf => N_428,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_388,
datab => \GRLFPC2_0.COMB.WRDATA_4\(22));
\GRLFPC2_0_COMB_WRDATA_4_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(32),
dataf => \GRLFPC2_0.R.I.RES\(29),
datae => \GRLFPC2_0.R.I.RES\(32),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(0),
dataf => N_406,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_366,
datab => \GRLFPC2_0.COMB.WRDATA_4\(32));
\GRLFPC2_0_COMB_WRDATA_4_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(34),
dataf => \GRLFPC2_0.R.I.RES\(31),
datae => \GRLFPC2_0.R.I.RES\(34),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(2),
dataf => N_408,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_368,
datab => \GRLFPC2_0.COMB.WRDATA_4\(34));
\GRLFPC2_0_COMB_WRDATA_4_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(36),
dataf => \GRLFPC2_0.R.I.RES\(33),
datae => \GRLFPC2_0.R.I.RES\(36),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(4),
dataf => N_410,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_370,
datab => \GRLFPC2_0.COMB.WRDATA_4\(36));
\GRLFPC2_0_COMB_DBGDATA_4_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(26),
dataf => \GRLFPC2_0.R.FSR.TEM\(3),
datae => N_400,
datad => N_401,
datac => N_692,
datab => N_628);
\GRLFPC2_0_COMB_WRDATA_4_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(5),
dataf => \GRLFPC2_0.R.I.RES\(34),
datae => \GRLFPC2_0.R.I.RES\(5),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(5),
dataf => N_411,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_371,
datab => \GRLFPC2_0.COMB.WRDATA_4\(5));
\GRLFPC2_0_COMB_WRDATA_4_14_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(14),
dataf => \GRLFPC2_0.R.I.RES\(43),
datae => \GRLFPC2_0.R.I.RES\(14),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_14_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(14),
dataf => N_420,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_380,
datab => \GRLFPC2_0.COMB.WRDATA_4\(14));
\GRLFPC2_0_COMB_WRDATA_4_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(17),
dataf => \GRLFPC2_0.R.I.RES\(46),
datae => \GRLFPC2_0.R.I.RES\(17),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(17),
dataf => N_423,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_383,
datab => \GRLFPC2_0.COMB.WRDATA_4\(17));
\GRLFPC2_0_COMB_WRDATA_4_20_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(20),
dataf => \GRLFPC2_0.R.I.RES\(49),
datae => \GRLFPC2_0.R.I.RES\(20),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_20_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(20),
dataf => N_426,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_386,
datab => \GRLFPC2_0.COMB.WRDATA_4\(20));
\GRLFPC2_0_COMB_WRDATA_4_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(24),
dataf => \GRLFPC2_0.R.I.RES\(53),
datae => \GRLFPC2_0.R.I.RES\(24),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(24),
dataf => N_430,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_390,
datab => \GRLFPC2_0.COMB.WRDATA_4\(24));
\GRLFPC2_0_COMB_WRDATA_4_37_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(37),
dataf => \GRLFPC2_0.R.I.RES\(34),
datae => \GRLFPC2_0.R.I.RES\(37),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_37_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(5),
dataf => N_411,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_371,
datab => \GRLFPC2_0.COMB.WRDATA_4\(37));
\GRLFPC2_0_COMB_WRDATA_4_46_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(46),
dataf => \GRLFPC2_0.R.I.RES\(43),
datae => \GRLFPC2_0.R.I.RES\(46),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_46_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(14),
dataf => N_420,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_380,
datab => \GRLFPC2_0.COMB.WRDATA_4\(46));
\GRLFPC2_0_COMB_WRDATA_4_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(49),
dataf => \GRLFPC2_0.R.I.RES\(46),
datae => \GRLFPC2_0.R.I.RES\(49),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(17),
dataf => N_423,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_383,
datab => \GRLFPC2_0.COMB.WRDATA_4\(49));
\GRLFPC2_0_COMB_WRDATA_4_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(52),
dataf => \GRLFPC2_0.R.I.RES\(49),
datae => \GRLFPC2_0.R.I.RES\(52),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(20),
dataf => N_426,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_386,
datab => \GRLFPC2_0.COMB.WRDATA_4\(52));
\GRLFPC2_0_COMB_WRDATA_4_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(56),
dataf => \GRLFPC2_0.R.I.RES\(53),
datae => \GRLFPC2_0.R.I.RES\(56),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(24),
dataf => N_430,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_390,
datab => \GRLFPC2_0.COMB.WRDATA_4\(56));
\GRLFPC2_0_COMB_DBGDATA_4_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(7),
dataf => \GRLFPC2_0.R.FSR.AEXC\(2),
datae => N_400,
datad => N_401,
datac => N_673,
datab => N_609);
\GRLFPC2_0_COMB_DBGDATA_4_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(25),
dataf => \GRLFPC2_0.R.FSR.TEM\(2),
datae => N_400,
datad => N_401,
datac => N_691,
datab => N_627);
\GRLFPC2_0_COMB_WRDATA_4_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(7),
dataf => \GRLFPC2_0.R.I.RES\(36),
datae => \GRLFPC2_0.R.I.RES\(7),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(7),
dataf => N_413,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_373,
datab => \GRLFPC2_0.COMB.WRDATA_4\(7));
\GRLFPC2_0_COMB_WRDATA_4_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(11),
dataf => \GRLFPC2_0.R.I.RES\(40),
datae => \GRLFPC2_0.R.I.RES\(11),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(11),
dataf => N_417,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_377,
datab => \GRLFPC2_0.COMB.WRDATA_4\(11));
\GRLFPC2_0_COMB_WRDATA_4_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(13),
dataf => \GRLFPC2_0.R.I.RES\(42),
datae => \GRLFPC2_0.R.I.RES\(13),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(13),
dataf => N_419,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_379,
datab => \GRLFPC2_0.COMB.WRDATA_4\(13));
\GRLFPC2_0_COMB_WRDATA_4_16_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(16),
dataf => \GRLFPC2_0.R.I.RES\(45),
datae => \GRLFPC2_0.R.I.RES\(16),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_16_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(16),
dataf => N_422,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_382,
datab => \GRLFPC2_0.COMB.WRDATA_4\(16));
\GRLFPC2_0_COMB_WRDATA_4_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(19),
dataf => \GRLFPC2_0.R.I.RES\(48),
datae => \GRLFPC2_0.R.I.RES\(19),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(19),
dataf => N_425,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_385,
datab => \GRLFPC2_0.COMB.WRDATA_4\(19));
\GRLFPC2_0_COMB_WRDATA_4_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(42),
dataf => \GRLFPC2_0.R.I.RES\(39),
datae => \GRLFPC2_0.R.I.RES\(42),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(10),
dataf => N_416,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_376,
datab => \GRLFPC2_0.COMB.WRDATA_4\(42));
\GRLFPC2_0_COMB_WRDATA_4_43_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(43),
dataf => \GRLFPC2_0.R.I.RES\(40),
datae => \GRLFPC2_0.R.I.RES\(43),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_43_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(11),
dataf => N_417,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_377,
datab => \GRLFPC2_0.COMB.WRDATA_4\(43));
\GRLFPC2_0_COMB_WRDATA_4_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(48),
dataf => \GRLFPC2_0.R.I.RES\(45),
datae => \GRLFPC2_0.R.I.RES\(48),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(16),
dataf => N_422,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_382,
datab => \GRLFPC2_0.COMB.WRDATA_4\(48));
\GRLFPC2_0_COMB_WRDATA_4_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(51),
dataf => \GRLFPC2_0.R.I.RES\(48),
datae => \GRLFPC2_0.R.I.RES\(51),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(19),
dataf => N_425,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_385,
datab => \GRLFPC2_0.COMB.WRDATA_4\(51));
\GRLFPC2_0_COMB_DBGDATA_4_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(1),
dataf => \GRLFPC2_0.R.FSR.CEXC\(1),
datae => N_400,
datad => N_401,
datac => N_667,
datab => N_603);
\GRLFPC2_0_COMB_DBGDATA_4_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(6),
dataf => \GRLFPC2_0.R.FSR.AEXC\(1),
datae => N_400,
datad => N_401,
datac => N_672,
datab => N_608);
\GRLFPC2_0_COMB_DBGDATA_4_30_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(30),
dataf => \GRLFPC2_0.R.FSR.RD\(0),
datae => N_400,
datad => N_401,
datac => N_696,
datab => N_632);
\GRLFPC2_0_COMB_WRDATA_4_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(6),
dataf => \GRLFPC2_0.R.I.RES\(35),
datae => \GRLFPC2_0.R.I.RES\(6),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(6),
dataf => N_412,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_372,
datab => \GRLFPC2_0.COMB.WRDATA_4\(6));
\GRLFPC2_0_COMB_WRDATA_4_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(12),
dataf => \GRLFPC2_0.R.I.RES\(41),
datae => \GRLFPC2_0.R.I.RES\(12),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(12),
dataf => N_418,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_378,
datab => \GRLFPC2_0.COMB.WRDATA_4\(12));
\GRLFPC2_0_COMB_WRDATA_4_30_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(30),
dataf => \GRLFPC2_0.R.I.RES\(59),
datae => \GRLFPC2_0.R.I.RES\(30),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_30_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(30),
dataf => N_436,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_396,
datab => \GRLFPC2_0.COMB.WRDATA_4\(30));
\GRLFPC2_0_COMB_WRDATA_4_35_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(35),
dataf => \GRLFPC2_0.R.I.RES\(32),
datae => \GRLFPC2_0.R.I.RES\(35),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_35_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(3),
dataf => N_409,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_369,
datab => \GRLFPC2_0.COMB.WRDATA_4\(35));
\GRLFPC2_0_COMB_WRDATA_4_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(38),
dataf => \GRLFPC2_0.R.I.RES\(35),
datae => \GRLFPC2_0.R.I.RES\(38),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(6),
dataf => N_412,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_372,
datab => \GRLFPC2_0.COMB.WRDATA_4\(38));
\GRLFPC2_0_COMB_WRDATA_4_44_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(44),
dataf => \GRLFPC2_0.R.I.RES\(41),
datae => \GRLFPC2_0.R.I.RES\(44),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_44_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(12),
dataf => N_418,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_378,
datab => \GRLFPC2_0.COMB.WRDATA_4\(44));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0ff00cccc")
port map (
combout => \GRLFPC2_0.N_3086\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.FSR.CEXC\(3),
datac => N_669,
datab => N_605);
\GRLFPC2_0_COMB_WRDATA_4_9_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(9),
dataf => \GRLFPC2_0.R.I.RES\(38),
datae => \GRLFPC2_0.R.I.RES\(9),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_9_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(9),
dataf => N_415,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_375,
datab => \GRLFPC2_0.COMB.WRDATA_4\(9));
\GRLFPC2_0_COMB_WRDATA_4_41_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(41),
dataf => \GRLFPC2_0.R.I.RES\(38),
datae => \GRLFPC2_0.R.I.RES\(41),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_41_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(9),
dataf => N_415,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_375,
datab => \GRLFPC2_0.COMB.WRDATA_4\(41));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcc3300fcfc3030")
port map (
combout => \GRLFPC2_0.N_3079\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.INST\(29),
datad => \GRLFPC2_0.FPCI_O\(312),
datac => \GRLFPC2_0.R.I.PC_O\(29),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_RS1_1_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => RFI2_RD1ADDRZ(0),
dataf => \GRLFPC2_0.COMB.RS1_1\(1),
datae => N_402,
datad => N_398);
\GRLFPC2_0_WRADDR_1_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRADDRZ(0),
dataf => N_402,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.WRADDR_1_SQMUXA\,
datac => \GRLFPC2_0.R.I.INST\(26),
datab => N_355);
\GRLFPC2_0_COMB_V_I_PC_1_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.R.I.PC\(25),
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.FPCI_O\(308),
datad => \GRLFPC2_0.R.I.PC_O\(25));
\GRLFPC2_0_COMB_V_I_PC_1_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.R.I.PC\(26),
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.FPCI_O\(309),
datad => \GRLFPC2_0.R.I.PC_O\(26));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_I_M2_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00fc30fc30")
port map (
combout => \GRLFPC2_0.N_3433\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.FPCI_O\(288),
datad => \GRLFPC2_0.R.I.INST\(5),
datac => \GRLFPC2_0.R.I.PC_O\(5),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_COMB_V_E_STDATA_1_0_I_M2_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00fc30fc30")
port map (
combout => \GRLFPC2_0.N_3434\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.FPCI_O\(294),
datad => \GRLFPC2_0.R.I.INST\(11),
datac => \GRLFPC2_0.R.I.PC_O\(11),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_COMB_V_E_STDATA_1_0_I_M2_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00fc30fc30")
port map (
combout => \GRLFPC2_0.N_3435\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.FPCI_O\(295),
datad => \GRLFPC2_0.R.I.INST\(12),
datac => \GRLFPC2_0.R.I.PC_O\(12),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_COMB_V_E_STDATA_1_0_I_M2_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00fc30fc30")
port map (
combout => \GRLFPC2_0.N_3436\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.FPCI_O\(296),
datad => \GRLFPC2_0.R.I.INST\(13),
datac => \GRLFPC2_0.R.I.PC_O\(13),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_COMB_V_E_STDATA_1_0_I_M2_15_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00fc30fc30")
port map (
combout => \GRLFPC2_0.N_3437\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.FPCI_O\(298),
datad => \GRLFPC2_0.R.I.INST\(15),
datac => \GRLFPC2_0.R.I.PC_O\(15),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_COMB_V_E_STDATA_1_0_I_M2_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00fc30fc30")
port map (
combout => \GRLFPC2_0.N_3439\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.FPCI_O\(300),
datad => \GRLFPC2_0.R.I.INST\(17),
datac => \GRLFPC2_0.R.I.PC_O\(17),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_COMB_V_I_PC_1_I_M2_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.N_3425\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.FPCI_O\(301),
datad => \GRLFPC2_0.R.I.PC_O\(18));
\GRLFPC2_0_COMB_V_I_PC_1_I_M2_20_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.N_3426\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.FPCI_O\(303),
datad => \GRLFPC2_0.R.I.PC_O\(20));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_I_M2_21_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00fc30fc30")
port map (
combout => \GRLFPC2_0.N_3442\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.FPCI_O\(304),
datad => \GRLFPC2_0.R.I.INST\(21),
datac => \GRLFPC2_0.R.I.PC_O\(21),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_COMB_V_E_STDATA_1_0_I_M2_22_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00fc30fc30")
port map (
combout => \GRLFPC2_0.N_3443\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.FPCI_O\(305),
datad => \GRLFPC2_0.R.I.INST\(22),
datac => \GRLFPC2_0.R.I.PC_O\(22),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_COMB_V_E_STDATA_1_0_I_M2_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00fc30fc30")
port map (
combout => \GRLFPC2_0.N_3445\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.FPCI_O\(307),
datad => \GRLFPC2_0.R.I.INST\(24),
datac => \GRLFPC2_0.R.I.PC_O\(24),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_COMB_V_E_STDATA_1_0_I_M2_30_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00fc30fc30")
port map (
combout => \GRLFPC2_0.N_3446\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.FPCI_O\(313),
datad => \GRLFPC2_0.R.I.INST\(30),
datac => \GRLFPC2_0.R.I.PC_O\(30),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_COMB_WRDATA_4_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(26),
dataf => \GRLFPC2_0.R.I.RES\(55),
datae => \GRLFPC2_0.R.I.RES\(26),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(26),
dataf => N_432,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_392,
datab => \GRLFPC2_0.COMB.WRDATA_4\(26));
\GRLFPC2_0_COMB_WRDATA_4_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(58),
dataf => \GRLFPC2_0.R.I.RES\(55),
datae => \GRLFPC2_0.R.I.RES\(58),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(26),
dataf => N_432,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_392,
datab => \GRLFPC2_0.COMB.WRDATA_4\(58));
\GRLFPC2_0_COMB_WRDATA_4_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(29),
dataf => \GRLFPC2_0.R.I.RES\(58),
datae => \GRLFPC2_0.R.I.RES\(29),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(29),
dataf => N_435,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_395,
datab => \GRLFPC2_0.COMB.WRDATA_4\(29));
\GRLFPC2_0_COMB_WRDATA_4_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(61),
dataf => \GRLFPC2_0.R.I.RES\(58),
datae => \GRLFPC2_0.R.I.RES\(61),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(29),
dataf => N_435,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_395,
datab => \GRLFPC2_0.COMB.WRDATA_4\(61));
\GRLFPC2_0_COMB_WRDATA_4_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(18),
dataf => \GRLFPC2_0.R.I.RES\(47),
datae => \GRLFPC2_0.R.I.RES\(18),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(18),
dataf => N_424,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_384,
datab => \GRLFPC2_0.COMB.WRDATA_4\(18));
\GRLFPC2_0_COMB_WRDATA_4_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(50),
dataf => \GRLFPC2_0.R.I.RES\(47),
datae => \GRLFPC2_0.R.I.RES\(50),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(18),
dataf => N_424,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_384,
datab => \GRLFPC2_0.COMB.WRDATA_4\(50));
\GRLFPC2_0_WRADDR_1_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRADDRZ(2),
dataf => N_404,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.WRADDR_1_SQMUXA\,
datac => \GRLFPC2_0.R.I.INST\(28),
datab => N_357);
\GRLFPC2_0_COMB_V_I_PC_1_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.R.I.PC\(3),
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.FPCI_O\(286),
datad => \GRLFPC2_0.R.I.PC_O\(3));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00fc30fc30")
port map (
combout => \GRLFPC2_0.N_3054\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.FPCI_O\(287),
datad => \GRLFPC2_0.R.I.INST\(4),
datac => \GRLFPC2_0.R.I.PC_O\(4),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_COMB_V_E_STDATA_1_0_9_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00fc30fc30")
port map (
combout => \GRLFPC2_0.N_3059\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.FPCI_O\(292),
datad => \GRLFPC2_0.R.I.INST\(9),
datac => \GRLFPC2_0.R.I.PC_O\(9),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_COMB_V_E_STDATA_1_0_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcc3300fcfc3030")
port map (
combout => \GRLFPC2_0.N_3069\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.INST\(19),
datad => \GRLFPC2_0.FPCI_O\(302),
datac => \GRLFPC2_0.R.I.PC_O\(19),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_COMB_DBGDATA_4_14_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(14),
dataf => \GRLFPC2_0.R.FSR.FTT\(0),
datae => N_400,
datad => N_401,
datac => N_680,
datab => N_616);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_RNIG14OGE3_68_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000f0f0f000f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0_N_5\,
dataf => N_27316,
datae => N_27258,
datad => N_27315,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIGJ2IDT2_0_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0_N_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0_M3_I_A3_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_RNIE3QJME3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"4c4c4c4444444c44")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_2\,
dataf => N_27316,
datae => N_27258,
datad => N_27315,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_112_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(112),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(112),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(112),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_111_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(111),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(111),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(111),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_110_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(110),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(110),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(110),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_107_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(107),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(107),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(107),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_106_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(106),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(106),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(106),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_103_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(103),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(103),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(103),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_101_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(101),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(101),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(101),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_93_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(93),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(93),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(93),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_91_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(91),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(91),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(91));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(83),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_82_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(82),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(82),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(82),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_81_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_78_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(78),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_75_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(75),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(75),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(75),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_73_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(73),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(73),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_70_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(70),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(70),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(70),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_69_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(69),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(69),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(69),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_68_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(68),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(68),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(68),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_67_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(67),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(67),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(67),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_66_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(66),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(66),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(66),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_65_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(65),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(65),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(65),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_63_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(63),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(63),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(63));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(62),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(62),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(62));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(61),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(61),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_113_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(113),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_112_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0ff00aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(112),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datad => \GRLFPC2_0.FPO.FRAC\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_111_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0ff00aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(111),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datad => \GRLFPC2_0.FPO.FRAC\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_110_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0ff00aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(110),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datad => \GRLFPC2_0.FPO.FRAC\(5),
datac => \GRLFPC2_0.FPO.FRAC\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_107_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0ff00aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(107),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datad => \GRLFPC2_0.FPO.FRAC\(8),
datac => \GRLFPC2_0.FPO.FRAC\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_106_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0ff00aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(106),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datad => \GRLFPC2_0.FPO.FRAC\(9),
datac => \GRLFPC2_0.FPO.FRAC\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_105_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(105),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datad => \GRLFPC2_0.FPO.FRAC\(10),
datac => \GRLFPC2_0.FPO.FRAC\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_104_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(104),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datad => \GRLFPC2_0.FPO.FRAC\(11),
datac => \GRLFPC2_0.FPO.FRAC\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_103_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0ff00aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(103),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datad => \GRLFPC2_0.FPO.FRAC\(12),
datac => \GRLFPC2_0.FPO.FRAC\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_102_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(102),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datad => \GRLFPC2_0.FPO.FRAC\(13),
datac => \GRLFPC2_0.FPO.FRAC\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_101_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0ff00aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(101),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datad => \GRLFPC2_0.FPO.FRAC\(14),
datac => \GRLFPC2_0.FPO.FRAC\(12),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_100_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(100),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datad => \GRLFPC2_0.FPO.FRAC\(15),
datac => \GRLFPC2_0.FPO.FRAC\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_99_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(99),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datad => \GRLFPC2_0.FPO.FRAC\(16),
datac => \GRLFPC2_0.FPO.FRAC\(14),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_98_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(98),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datad => \GRLFPC2_0.FPO.FRAC\(17),
datac => \GRLFPC2_0.FPO.FRAC\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_97_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(97),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datad => \GRLFPC2_0.FPO.FRAC\(18),
datac => \GRLFPC2_0.FPO.FRAC\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_94_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(94),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datad => \GRLFPC2_0.FPO.FRAC\(21),
datac => \GRLFPC2_0.FPO.FRAC\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_93_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0ff00aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(93),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datad => \GRLFPC2_0.FPO.FRAC\(22),
datac => \GRLFPC2_0.FPO.FRAC\(20),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_92_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(92),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datad => \GRLFPC2_0.FPO.FRAC\(23),
datac => \GRLFPC2_0.FPO.FRAC\(21),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_91_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0ff00aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(91),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datad => \GRLFPC2_0.FPO.FRAC\(24),
datac => \GRLFPC2_0.FPO.FRAC\(22),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_90_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(90),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datad => \GRLFPC2_0.FPO.FRAC\(25),
datac => \GRLFPC2_0.FPO.FRAC\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_89_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(89),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datad => \GRLFPC2_0.FPO.FRAC\(26),
datac => \GRLFPC2_0.FPO.FRAC\(24),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_88_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(88),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datad => \GRLFPC2_0.FPO.FRAC\(27),
datac => \GRLFPC2_0.FPO.FRAC\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_87_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(87),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datad => \GRLFPC2_0.FPO.FRAC\(28),
datac => \GRLFPC2_0.FPO.FRAC\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_86_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(86),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datad => \GRLFPC2_0.FPO.FRAC\(29),
datac => \GRLFPC2_0.FPO.FRAC\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_85_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaff00f0f0cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(85),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(30),
datac => \GRLFPC2_0.FPO.FRAC\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_84_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaff00f0f0cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(84),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(31),
datac => \GRLFPC2_0.FPO.FRAC\(29),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccff00f0f0aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(83),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(30),
datac => \GRLFPC2_0.FPO.FRAC\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_82_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(82),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(33),
datac => \GRLFPC2_0.FPO.FRAC\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_81_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0ff00aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(34),
datac => \GRLFPC2_0.FPO.FRAC\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_79_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(36),
datac => \GRLFPC2_0.FPO.FRAC\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_78_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0ff00aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(78),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(37),
datac => \GRLFPC2_0.FPO.FRAC\(35),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_77_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(77),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(38),
datac => \GRLFPC2_0.FPO.FRAC\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_76_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(76),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(39),
datac => \GRLFPC2_0.FPO.FRAC\(37),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_75_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0ff00aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(75),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(40),
datac => \GRLFPC2_0.FPO.FRAC\(38),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_74_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(74),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(41),
datac => \GRLFPC2_0.FPO.FRAC\(39),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_73_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccff00f0f0aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(73),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(40),
datac => \GRLFPC2_0.FPO.FRAC\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_70_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(70),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(45),
datac => \GRLFPC2_0.FPO.FRAC\(43),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_69_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(69),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(46),
datac => \GRLFPC2_0.FPO.FRAC\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_68_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0ff00aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(68),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(47),
datac => \GRLFPC2_0.FPO.FRAC\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_67_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0ff00aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(67),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(48),
datac => \GRLFPC2_0.FPO.FRAC\(46),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_66_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0ff00aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(66),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(49),
datac => \GRLFPC2_0.FPO.FRAC\(47),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_65_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0ff00aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(65),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(50),
datac => \GRLFPC2_0.FPO.FRAC\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_63_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0ff00aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(63),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(52),
datac => \GRLFPC2_0.FPO.FRAC\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0ff00aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(62),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(53),
datac => \GRLFPC2_0.FPO.FRAC\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0ff00aaaa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(61),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(54),
datac => \GRLFPC2_0.FPO.FRAC\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_114_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000c000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(114),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(117));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIU3R3OL_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(29),
dataf => N_27258,
datae => N_27260,
datad => N_27259);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIM296PL_30_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(30),
dataf => N_27258,
datae => N_27261,
datad => N_27262);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIK6L6RL_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(31),
dataf => N_27258,
datae => N_27264,
datad => N_27263);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIKED7VL_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(32),
dataf => N_27258,
datae => N_27266,
datad => N_27265);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI4VUBNM_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(34),
dataf => N_27258,
datae => N_27270,
datad => N_27269);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIS15UNP_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(36),
dataf => N_27258,
datae => N_27274,
datad => N_27273);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIO5DMOT_37_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(37),
dataf => N_27258,
datae => N_27276,
datad => N_27275);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIGCV93M2_40_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(40),
dataf => N_27258,
datae => N_27282,
datad => N_27281);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIKA2EFM_41_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(41),
dataf => N_27258,
datae => N_27284,
datad => N_27283);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI078M7N_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(42),
dataf => N_27258,
datae => N_27286,
datad => N_27285);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNISVJ6OO_43_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(43),
dataf => N_27258,
datae => N_27288,
datad => N_27287);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIOHB7PR_44_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(44),
dataf => N_27258,
datae => N_27290,
datad => N_27289);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIEO2SU11_45_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(45),
dataf => N_27258,
datae => N_27292,
datad => N_27291);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI439I6E1_46_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(46),
dataf => N_27258,
datae => N_27294,
datad => N_27293);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_15: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_15\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_22: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000300000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_22\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_15\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_26: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0003000f00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_26\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_22\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_20: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_20\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_19: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_19\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_17: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_17\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_23: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000300000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_23\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_17\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_27: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0003000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_27\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_23\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_19\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_252_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfffcf00c0ffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10522\,
dataf => \GRLFPC2_0.FPO.EXP\(6),
datae => \GRLFPC2_0.FPO.EXP\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(239));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_251_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfffcf00c0ffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10523\,
dataf => \GRLFPC2_0.FPO.EXP\(7),
datae => \GRLFPC2_0.FPO.EXP\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(238));
\GRLFPC2_0_COMB_DBGDATA_4_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff00f0f0")
port map (
combout => CPO_DBG_DATAZ(19),
dataf => N_400,
datae => N_401,
datad => N_685,
datac => N_621);
\GRLFPC2_0_COMB_DBGDATA_4_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff00f0f0")
port map (
combout => CPO_DBG_DATAZ(28),
dataf => N_400,
datae => N_401,
datad => N_694,
datac => N_630);
\GRLFPC2_0_COMB_V_E_STDATA_1_0_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33cc00fc30fc30")
port map (
combout => \GRLFPC2_0.N_3052\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.FPCI_O\(285),
datad => \GRLFPC2_0.R.I.INST\(2),
datac => \GRLFPC2_0.R.I.PC_O\(2),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_COMB_V_I_PC_1_I_M2_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.N_3432\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.FPCI_O\(314),
datad => \GRLFPC2_0.R.I.PC_O\(31));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0ff00cccc")
port map (
combout => \GRLFPC2_0.N_3114\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.FSR.RD\(1),
datac => N_697,
datab => N_633);
\GRLFPC2_0_COMB_DBGDATA_4_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(31),
dataf => \GRLFPC2_0.R.FSR.RD\(1),
datae => N_400,
datad => N_401,
datac => N_697,
datab => N_633);
\GRLFPC2_0_COMB_DBGDATA_4_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(2),
dataf => \GRLFPC2_0.R.FSR.CEXC\(2),
datae => N_400,
datad => N_401,
datac => N_668,
datab => N_604);
GRLFPC2_0_V_FSR_CEXC_3_SQMUXA: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000000f")
port map (
combout => \GRLFPC2_0.V.FSR.CEXC_3_SQMUXA\,
dataf => \GRLFPC2_0.N_1439\,
datae => \GRLFPC2_0.N_1015\,
datad => \GRLFPC2_0.N_1171\,
datac => \GRLFPC2_0.N_1517\);
GRLFPC2_0_R_I_V_ENA_RNO_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff00ff")
port map (
combout => \GRLFPC2_0.R.I.V_1_0_G0_I_O4_1\,
dataf => \GRLFPC2_0.N_1015\,
datae => \GRLFPC2_0.COMB.ANNULRES_1\,
datad => N_11);
GRLFPC2_0_COMB_ANNULRES_1_IV: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3f0c3f0f3f0c3300")
port map (
combout => \GRLFPC2_0.COMB.ANNULRES_1\,
dataf => \GRLFPC2_0.N_82\,
datae => \GRLFPC2_0.R.X.FPOP\,
datad => \GRLFPC2_0.R.X.SEQERR\,
datac => \GRLFPC2_0.R.I.EXEC\,
datab => \GRLFPC2_0.N_1105\);
GRLFPC2_0_R_I_V_ENA: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ff00fc0c")
port map (
combout => N_38488,
dataf => \GRLFPC2_0.N_1439\,
datae => \GRLFPC2_0.N_1876_2\,
datad => \GRLFPC2_0.R.I.V_1_0_G2\,
datac => \GRLFPC2_0.R.I.V_1_0_G0_I_O4_1\,
datab => \GRLFPC2_0.R.I.V\);
\GRLFPC2_0_WRDATA_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(1),
dataf => N_407,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_367,
datab => \GRLFPC2_0.COMB.WRDATA_4\(33));
\GRLFPC2_0_WRDATA_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(1),
dataf => N_407,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_367,
datab => \GRLFPC2_0.COMB.WRDATA_4\(1));
\GRLFPC2_0_COMB_WRDATA_4_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(33),
dataf => \GRLFPC2_0.R.I.RES\(30),
datae => \GRLFPC2_0.R.I.RES\(33),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_COMB_WRDATA_4_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(1),
dataf => \GRLFPC2_0.R.I.RES\(30),
datae => \GRLFPC2_0.R.I.RES\(1),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(4),
dataf => N_410,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_370,
datab => \GRLFPC2_0.COMB.WRDATA_4\(4));
\GRLFPC2_0_COMB_WRDATA_4_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(4),
dataf => \GRLFPC2_0.R.I.RES\(33),
datae => \GRLFPC2_0.R.I.RES\(4),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_COMB_RS2_1_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000fffff0000000")
port map (
combout => \GRLFPC2_0.COMB.RS2_1\(1),
dataf => \GRLFPC2_0.R.A.RS2\(1),
datae => N_13,
datad => \GRLFPC2_0.N_951\,
datac => N_54);
GRLFPC2_0_COMB_UN1_MEXC_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f00ff0f0fffff")
port map (
combout => \GRLFPC2_0.COMB.UN1_MEXC_0\,
dataf => \GRLFPC2_0.R.FSR.TEM\(0),
datae => \GRLFPC2_0.R.FSR.TEM\(3),
datad => \GRLFPC2_0.R.I.EXC\(0),
datac => \GRLFPC2_0.R.I.EXC\(3));
GRLFPC2_0_COMB_UN1_MEXC_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f00ff0f0fffff")
port map (
combout => \GRLFPC2_0.COMB.UN1_MEXC_1\,
dataf => \GRLFPC2_0.R.FSR.TEM\(1),
datae => \GRLFPC2_0.R.FSR.TEM\(4),
datad => \GRLFPC2_0.R.I.EXC\(1),
datac => \GRLFPC2_0.R.I.EXC\(4));
GRLFPC2_0_R_I_EXEC_RNO_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000ff00ff00ff00")
port map (
combout => N_37320,
dataf => \GRLFPC2_0.COMB.UN1_MEXC_1\,
datae => \GRLFPC2_0.COMB.UN1_MEXC_0\,
datad => \GRLFPC2_0.R.I.V\,
datac => \GRLFPC2_0.R.FSR.TEM\(2),
datab => \GRLFPC2_0.R.I.EXC\(2));
GRLFPC2_0_COMB_V_I_RDD_1_I_A3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.N_1438\,
dataf => \GRLFPC2_0.N_1438_15\,
datae => N_13);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"5050f0005353f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIG3MJ_40_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4662\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(39),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(40));
\GRLFPC2_0_WRDATA_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(28),
dataf => N_434,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_394,
datab => \GRLFPC2_0.COMB.WRDATA_4\(60));
\GRLFPC2_0_WRDATA_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(25),
dataf => N_431,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_391,
datab => \GRLFPC2_0.COMB.WRDATA_4\(57));
\GRLFPC2_0_WRDATA_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(28),
dataf => N_434,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_394,
datab => \GRLFPC2_0.COMB.WRDATA_4\(28));
\GRLFPC2_0_WRDATA_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRDATAZ(25),
dataf => N_431,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_391,
datab => \GRLFPC2_0.COMB.WRDATA_4\(25));
\GRLFPC2_0_COMB_WRDATA_4_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(60),
dataf => \GRLFPC2_0.R.I.RES\(57),
datae => \GRLFPC2_0.R.I.RES\(60),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_COMB_WRDATA_4_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(57),
dataf => \GRLFPC2_0.R.I.RES\(54),
datae => \GRLFPC2_0.R.I.RES\(57),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_COMB_WRDATA_4_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(28),
dataf => \GRLFPC2_0.R.I.RES\(57),
datae => \GRLFPC2_0.R.I.RES\(28),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_COMB_WRDATA_4_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(25),
dataf => \GRLFPC2_0.R.I.RES\(54),
datae => \GRLFPC2_0.R.I.RES\(25),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_WRDATA_45_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(13),
dataf => N_419,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_379,
datab => \GRLFPC2_0.COMB.WRDATA_4\(45));
\GRLFPC2_0_WRDATA_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI1_WRDATAZ(7),
dataf => N_413,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.N_1243\,
datac => N_373,
datab => \GRLFPC2_0.COMB.WRDATA_4\(39));
\GRLFPC2_0_COMB_WRDATA_4_45_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(45),
dataf => \GRLFPC2_0.R.I.RES\(42),
datae => \GRLFPC2_0.R.I.RES\(45),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_COMB_WRDATA_4_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4\(39),
dataf => \GRLFPC2_0.R.I.RES\(36),
datae => \GRLFPC2_0.R.I.RES\(39),
datad => \GRLFPC2_0.N_83\);
\GRLFPC2_0_COMB_DBGDATA_4_1_M3_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(13),
dataf => \GRLFPC2_0.N_76_I\,
datae => N_400,
datad => N_401,
datac => N_679,
datab => N_615);
\GRLFPC2_0_COMB_RF1REN_1_0_0_A2_1_0_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000f000000000")
port map (
combout => \GRLFPC2_0.N_77_1\,
dataf => \GRLFPC2_0.N_44\,
datae => N_66,
datad => N_58,
datac => N_59);
\GRLFPC2_0_COMB_V_A_RF2REN_1_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f000f000f0000")
port map (
combout => \GRLFPC2_0.COMB.V.A.RF2REN_1\(1),
dataf => \GRLFPC2_0.COMB.RS1D_1\,
datae => \GRLFPC2_0.COMB.RS1_1\(0),
datad => \GRLFPC2_0.N_3477_1_I\,
datac => N_37362);
\GRLFPC2_0_COMB_V_A_RF1REN_1_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f000f0000000f")
port map (
combout => \GRLFPC2_0.COMB.V.A.RF1REN_1\(1),
dataf => \GRLFPC2_0.COMB.RS1D_1\,
datae => \GRLFPC2_0.COMB.RS1_1\(0),
datad => \GRLFPC2_0.N_3477_1_I\,
datac => N_37362);
GRLFPC2_0_COMB_RS2D_1_IV_0_O2_RNII95D: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000c000000")
port map (
combout => \GRLFPC2_0.COMB.RS2D_1\,
dataf => N_66,
datae => \GRLFPC2_0.N_951\,
datad => \GRLFPC2_0.N_44\,
datac => N_58,
datab => N_59);
\GRLFPC2_0_COMB_RS2_1_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000fffff0000000")
port map (
combout => \GRLFPC2_0.COMB.RS2_1\(0),
dataf => \GRLFPC2_0.R.A.RS2\(0),
datae => N_13,
datad => \GRLFPC2_0.N_951\,
datac => N_53);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(58),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_176__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIOUT87M_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(33),
dataf => N_27258,
datae => N_27268,
datad => N_27267);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI001INN_35_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(35),
dataf => N_27258,
datae => N_27272,
datad => N_27271);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_80_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(35),
datac => \GRLFPC2_0.FPO.FRAC\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_96_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(96),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datad => \GRLFPC2_0.FPO.FRAC\(19),
datac => \GRLFPC2_0.FPO.FRAC\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf3f0ff0c03000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(2),
datae => N_53980,
datad => N_53982,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"333ff3ff000cc0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(56),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f0ff00ff00")
port map (
combout => N_53942,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff0ffff0ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_O2_1_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0fff0f0cffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN11_WQSTSETS\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00fff0ff0fffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(56),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8_I\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00fff0ff0fffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_95_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaf0f0ff00cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(95),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0\,
datad => \GRLFPC2_0.FPO.FRAC\(20),
datac => \GRLFPC2_0.FPO.FRAC\(18),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53882,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbcbf8c83b0b3808")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10038\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(36),
datae => \GRLFPC2_0.FPO.FRAC\(21),
datad => \GRLFPC2_0.FPO.FRAC\(20),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_247_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfffc0ffcf00c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10527\,
dataf => \GRLFPC2_0.FPO.EXP\(10),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_249_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfffcf00c0ffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10525\,
dataf => \GRLFPC2_0.FPO.EXP\(9),
datae => \GRLFPC2_0.FPO.EXP\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3639\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_CIN_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33f0cc00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6583\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_58_0_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cf3fffff30c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58\(56),
dataf => N_30731,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5771\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_0_RNIIUSV: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff00ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1281_I\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1274_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_CIN_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33f0cc00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5771\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_CIN_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33f0cc00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6583\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_SA_I_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cf3f30cffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1_0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fccf000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5771\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(57),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(316));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"330fccf000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10626\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(258));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_0_RNIIUSV_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0000ff00ffff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.56.SI_60\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1274_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_55_CI_60_Z_1_CO1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffccc0fcc0fccc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_60.Z_1_CO1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1274_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN_2\);
GRLFPC2_0_R_A_FPOP_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000c0f00000c0c0")
port map (
combout => \GRLFPC2_0.R.A.FPOP_0_0_G1\,
dataf => \GRLFPC2_0.N_1714_I\,
datae => \GRLFPC2_0.N_67\,
datad => \GRLFPC2_0.N_1093\,
datac => \GRLFPC2_0.N_951\,
datab => \GRLFPC2_0.N_1072\);
GRLFPC2_0_FPI_LDOP_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000ffff")
port map (
combout => \GRLFPC2_0.FPI.RST_1\,
dataf => \GRLFPC2_0.R.MK.RST2\,
datae => N_11);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_232__G2_0_7920_I_A7_7\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7920_I_A7_7\,
dataf => \GRLFPC2_0.FPCI_O_3\(74),
datae => \GRLFPC2_0.FPCI_O_0\(60),
datad => \GRLFPC2_0.FPCI_O_0\(69),
datac => \GRLFPC2_0.FPCI_O_0\(70));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_232__G2_0_7920_I_A7_10\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7920_I_A7_10\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7920_I_A7_7\,
datae => \GRLFPC2_0.HOLDN_O\,
datad => \GRLFPC2_0.FPCI_O_0\(61),
datac => \GRLFPC2_0.FPCI_O_0\(62),
datab => \GRLFPC2_0.FPCI_O_0\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_232__G2_0_7920_I_A7_6\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7920_I_A7_6\,
dataf => \GRLFPC2_0.FPCI_O_3\(0),
datae => \GRLFPC2_0.FPCI_O_0\(63),
datad => \GRLFPC2_0.FPCI_O_3\(73),
datac => \GRLFPC2_0.COMB.LOCKGEN.LOCKI_O_3\);
GRLFPC2_0_FPI_LDOP_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff3000000")
port map (
combout => \GRLFPC2_0.FPI.LDOP_1\,
dataf => \GRLFPC2_0.R.MK.RST\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7920_I_A7_10\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7920_I_A7_6\,
datac => \GRLFPC2_0.R.STATE_O_3\(1),
datab => \GRLFPC2_0.R.STATE_O_3\(0));
GRLFPC2_0_R_MK_HOLDN1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffffffff")
port map (
combout => \GRLFPC2_0.N_2103\,
dataf => \GRLFPC2_0.R.MK.RST2\,
datae => N_11);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_37_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000f030f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1496\,
dataf => N_28511,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_I_O2_3_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_118_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_33_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffc00000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1836\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_429\,
datad => N_35133,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_30_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000fffffff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1771\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_O2_14_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffc0ffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1844\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
datae => N_35133,
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_38_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffc000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1497\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_875\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_65_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fffcfffcfffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1495\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_875\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN2_DIVMULTV_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000f0000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_DIVMULTV\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_GRFPUF_0_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffcff00003000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(2),
dataf => \GRLFPC2_0.FPO.FRAC\(53),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_2_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00fc30ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_GRFPUF_0_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffcff00003000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(3),
dataf => \GRLFPC2_0.FPO.FRAC\(52),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_GRFPUF_0_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffcff00003000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(1),
dataf => \GRLFPC2_0.FPO.FRAC\(54),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_GRFPUF_0_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000300ffffcfff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_176__G2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_2_RNITA48_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000f0cc0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(375),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SIGNRESULT: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cccc0003c3cc0c")
port map (
combout => \GRLFPC2_0.FPO.SIGN\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(24),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_2_IV_1_TZ_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03030300cfcfcfcc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_IV_1_TZ\(0),
dataf => \GRLFPC2_0.FPO.SIGN\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4238\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNI1H4D_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4238\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_RNI9UPKME3_68_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0f0303030f030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4534\,
dataf => N_27316,
datae => N_27258,
datad => N_27315,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_2_IV_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00005a3300005aff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_I_I_0\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4534\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_I_M\(12),
datad => \GRLFPC2_0.FPI.LDOP_0\,
datac => \GRLFPC2_0.FPI.OP2\(63),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_IV_1_TZ\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f00088880f004444")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4874\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_I_I_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP\,
datad => N_36986,
datac => N_36985,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN53_SCTRL_NEW: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff03030303")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP\,
datae => N_36986,
datad => N_36985,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNI8T8G_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff0fffffff00")
port map (
combout => N_36986,
dataf => \GRLFPC2_0.R.FSR.RD\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(21),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN17_U_RDN_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff00")
port map (
combout => N_36985,
dataf => \GRLFPC2_0.R.FSR.RD\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(21),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI4NDI_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03300cc0300cc003")
port map (
combout => N_53997,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN2_MIXOIN_RNID1AV1_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00033cc03cc00003")
port map (
combout => N_53999,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SALSBS_1\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP_1_1_CO1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SALSBS_2\(0),
datac => N_53996,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5446\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN36_STKGEN_0_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00000000ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN36_STKGEN_0_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SCLSBS_1\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_954\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(373));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN2_MIXOIN_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcfcccccc0c000")
port map (
combout => N_53996,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN2_MIXOIN_1_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffcc0fcc00000")
port map (
combout => N_53998,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SALSBS_1\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP_1_1_CO1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SALSBS_2\(0),
datac => N_53996,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5446\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN2_MIXOIN_2_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffcc0fcc00000")
port map (
combout => N_54002,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SBLSBS_1\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_959_I\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SBLSBS_2\(0),
datac => N_53998,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5452\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN2_MIXOIN_3_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"edede848ffffa000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_3_I\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN25_NOTPROP\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_CARRY_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN26_GEN\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SCLSBS_2\(0),
datab => N_54002,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5458\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI3UVA_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cf3f30cf30cf30c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SALSBS_1\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(369));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIQOLG_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0c0c000c000c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP_1_1_CO1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(370));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00fff0f00000f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(312));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIQOLG_0_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cf3f30cf30cf30c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SALSBS_2\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(370));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(371));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f000f0fff000f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(313));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f000f0fff000f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(314));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN26_GEN: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN26_GEN\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SCLSBS_1\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_954\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00fff0f00000f0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(311));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI3UVA_0_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0c0c000c000c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_1_CO0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(369));
GRLFPC2_0_RS2_0_SQMUXA_0_0_A2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff000000")
port map (
combout => \GRLFPC2_0.N_3462\,
dataf => N_75,
datae => N_84,
datad => N_77);
GRLFPC2_0_UN1_FPOP7_1_0_A2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c00000000000000")
port map (
combout => \GRLFPC2_0.N_74\,
dataf => \GRLFPC2_0.N_3468\,
datae => \GRLFPC2_0.N_3466\,
datad => \GRLFPC2_0.N_951\,
datac => N_59,
datab => N_58);
GRLFPC2_0_UN1_FPOP7_1_0_A2_0_4: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000c0000000")
port map (
combout => \GRLFPC2_0.UN1_FPOP7_1_0_A2_0_2\,
dataf => N_60,
datae => N_61,
datad => \GRLFPC2_0.N_3468\,
datac => N_64,
datab => N_58);
GRLFPC2_0_UN1_FPOP7_1_0_A2_0_4_RNI1MSO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cfcfcf00ffffff")
port map (
combout => \GRLFPC2_0.COMB.V.A.RF1REN_1_8000_I_A5_0\,
dataf => \GRLFPC2_0.UN1_FPOP7_1_0_A2_0_2\,
datae => \GRLFPC2_0.RS1V_0_SQMUXA\,
datad => \GRLFPC2_0.N_1072\,
datac => \GRLFPC2_0.N_951\,
datab => N_59);
GRLFPC2_0_UN1_FPOP7_1_0_A2_RNILOL71: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000fff00000000")
port map (
combout => N_37362,
dataf => \GRLFPC2_0.COMB.V.A.RF1REN_1_8000_I_A5_0\,
datae => \GRLFPC2_0.N_74\,
datad => \GRLFPC2_0.N_951\,
datac => N_72);
GRLFPC2_0_COMB_FPDECODE_RS1D5_0_A2_0_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000c000000000000")
port map (
combout => \GRLFPC2_0.COMB.FPDECODE.RS1D5_0_A2_0\,
dataf => \GRLFPC2_0.N_3466\,
datae => N_62,
datad => N_66,
datac => N_58,
datab => N_59);
GRLFPC2_0_COMB_RS1D_1_U: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3f3f3fc0000000")
port map (
combout => \GRLFPC2_0.COMB.RS1D_1\,
dataf => \GRLFPC2_0.RS1D_CNST\,
datae => \GRLFPC2_0.COMB.FPDECODE.RS1D5_1\,
datad => \GRLFPC2_0.COMB.FPDECODE.RS1D5_0_A2_0\,
datac => \GRLFPC2_0.N_951\,
datab => N_72);
\GRLFPC2_0_COMB_RS1_1_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcfcfcf30000000")
port map (
combout => \GRLFPC2_0.COMB.RS1_1\(0),
dataf => \GRLFPC2_0.N_2975\,
datae => \GRLFPC2_0.RS1V_0_SQMUXA\,
datad => N_78,
datac => N_13,
datab => \GRLFPC2_0.N_951\);
GRLFPC2_0_RS1V_0_SQMUXA: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300000000000000")
port map (
combout => \GRLFPC2_0.RS1V_0_SQMUXA\,
dataf => N_84,
datae => N_83,
datad => \GRLFPC2_0.RS1V12_TZ\,
datac => N_76,
datab => N_75);
\GRLFPC2_0_R_A_RF1REN_RNO_0_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff000000")
port map (
combout => N_37365_1,
dataf => \GRLFPC2_0.RS1D_CNST\,
datae => \GRLFPC2_0.RS1V_0_SQMUXA\,
datad => N_78);
\GRLFPC2_0_COMB_RS1_1_0_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.N_2975\,
dataf => \GRLFPC2_0.R.A.RS1\(0),
datae => N_67,
datad => N_13);
GRLFPC2_0_COMB_RDD_1_M7_E_54_I_A2_0_4: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000ff00000000000")
port map (
combout => \GRLFPC2_0.COMB.RDD_1.M7_E_54_I_A2_0\,
dataf => \GRLFPC2_0.N_3468\,
datae => N_59,
datad => N_64,
datac => N_58);
GRLFPC2_0_COMB_RDD_1_M7_E_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f3ffffff")
port map (
combout => \GRLFPC2_0.COMB.RDD_1.M7_E_0\,
dataf => \GRLFPC2_0.N_925\,
datae => \GRLFPC2_0.COMB.RDD_1.M7_E_54_I_A2_0\,
datad => N_63,
datac => N_60,
datab => N_61);
GRLFPC2_0_COMB_RDD_1_M7_E_54_I_A2_0_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000f0000")
port map (
combout => \GRLFPC2_0.COMB.RDD_1.M7_E_54_I_A2_0_3\,
dataf => N_62,
datae => N_65,
datad => N_66,
datac => N_59);
GRLFPC2_0_COMB_RDD_1_M7_E: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3ffffff00000000")
port map (
combout => \GRLFPC2_0.COMB.RDD_1.N_27\,
dataf => \GRLFPC2_0.COMB.RDD_1.M7_E_0\,
datae => \GRLFPC2_0.COMB.RDD_1.M7_E_54_I_A2_0_3\,
datad => \GRLFPC2_0.N_3466\,
datac => N_60,
datab => N_61);
GRLFPC2_0_COMB_FPDECODE_RS1D5_0_A2_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => \GRLFPC2_0.COMB.FPDECODE.RS1D5_1\,
dataf => N_61,
datae => N_65);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_MIFROMINST_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f03030f0003030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.MIFROMINST_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(71),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(74));
GRLFPC2_0_COMB_V_MK_RST_1_4: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000000000000000")
port map (
combout => \GRLFPC2_0.R.MK.RST_4\,
dataf => \GRLFPC2_0.R.MK.HOLDN2\,
datae => \GRLFPC2_0.HOLDN_O\,
datad => \GRLFPC2_0.FPO.BUSY_O\,
datac => \GRLFPC2_0.R.MK.HOLDN2_O\);
GRLFPC2_0_COMB_V_MK_RST_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000f000000000")
port map (
combout => \GRLFPC2_0.R.MK.RST\,
dataf => \GRLFPC2_0.R.MK.RST_4\,
datae => \GRLFPC2_0.R.MK.RST2\,
datad => \GRLFPC2_0.R.MK.RST2_O\,
datac => \GRLFPC2_0.COMB.ANNULFPU_1_O\);
GRLFPC2_0_COMB_RSDECODE_RS1V: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => \GRLFPC2_0.N_1072\,
dataf => N_85,
datae => N_86);
GRLFPC2_0_COMB_LOCKGEN_UN8_DEPCHECK: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff0")
port map (
combout => \GRLFPC2_0.N_1093\,
dataf => \GRLFPC2_0.R.X.LD\,
datae => \GRLFPC2_0.R.A.LD\,
datad => \GRLFPC2_0.R.M.LD\,
datac => \GRLFPC2_0.R.E.LD\);
\GRLFPC2_0_COMB_RF1REN_1_0_0_A2_2_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000f000c000c000")
port map (
combout => \GRLFPC2_0.N_3475\,
dataf => \GRLFPC2_0.N_1714_I\,
datae => \GRLFPC2_0.N_1093\,
datad => N_13,
datac => \GRLFPC2_0.N_951\,
datab => \GRLFPC2_0.N_1072\);
GRLFPC2_0_FPI_START_0_A2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f00000000")
port map (
combout => \GRLFPC2_0.FPI.START\,
dataf => \GRLFPC2_0.N_3475\,
datae => \GRLFPC2_0.R.MK.RST\,
datad => \GRLFPC2_0.N_67\,
datac => \GRLFPC2_0.R.MK.RST2\);
GRLFPC2_0_RS1D_CNST_0_A2_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.N_624_3\,
dataf => N_74,
datae => N_77);
GRLFPC2_0_RS1D_CNST_0_A2_2_RNI8PIU: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000c000")
port map (
combout => \GRLFPC2_0.COMB.FPDECODE.ST\,
dataf => N_76,
datae => N_75,
datad => \GRLFPC2_0.N_624_3\,
datac => N_84,
datab => N_83);
GRLFPC2_0_COMB_FPDECODE_LD_0_O2_I_O2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000ffff")
port map (
combout => \GRLFPC2_0.N_45\,
dataf => N_72,
datae => N_73);
GRLFPC2_0_COMB_RS2D_1_IV_0_O2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff000000ff303030")
port map (
combout => \GRLFPC2_0.N_44\,
dataf => N_72,
datae => \GRLFPC2_0.N_3466\,
datad => \GRLFPC2_0.N_43\,
datac => \GRLFPC2_0.N_40\,
datab => N_60);
GRLFPC2_0_COMB_RS2D_1_IV_0_O2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000c30000000")
port map (
combout => \GRLFPC2_0.N_40\,
dataf => N_61,
datae => N_65,
datad => N_62,
datac => N_64,
datab => N_63);
GRLFPC2_0_COMB_RS2D_1_IV_0_O2_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000f0000f0c0f")
port map (
combout => \GRLFPC2_0.N_43\,
dataf => N_72,
datae => N_61,
datad => N_65,
datac => N_62,
datab => N_60);
GRLFPC2_0_UN1_FPOP7_1_0_A2_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000ff")
port map (
combout => \GRLFPC2_0.N_3468\,
dataf => N_66,
datae => N_65,
datad => N_62);
GRLFPC2_0_COMB_FPDECODE_RS1D5_0_A2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => \GRLFPC2_0.N_3466\,
dataf => N_64,
datae => N_63);
GRLFPC2_0_RS1D_CNST_0_O2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f0000c000c000")
port map (
combout => \GRLFPC2_0.N_2888\,
dataf => N_76,
datae => \GRLFPC2_0.N_925\,
datad => N_83,
datac => N_73,
datab => N_72);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MAPMULXFF_UN4_UNIMPMAP: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ffffffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7226\,
dataf => N_64,
datae => N_62,
datad => N_65);
GRLFPC2_0_COMB_PEXC8_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => CPO_EXCZ,
dataf => \GRLFPC2_0.R.STATE\(0),
datae => \GRLFPC2_0.R.STATE\(1));
\GRLFPC2_0_COMB_V_STATE_1_IV_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0c0f00000c00000")
port map (
combout => \GRLFPC2_0.R.STATE_0_0_1__I0_I_1\,
dataf => \GRLFPC2_0.N_1495\,
datae => \GRLFPC2_0.R.STATE\(0),
datad => \GRLFPC2_0.R.STATE\(1),
datac => \GRLFPC2_0.N_1667\,
datab => N_15);
GRLFPC2_0_COMB_V_I_RDD_1_I_A3_15_9: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000f000")
port map (
combout => \GRLFPC2_0.COMB.V.I.RDD_1_I_A3_15_9\,
dataf => \GRLFPC2_0.FPCI_O\(58),
datae => \GRLFPC2_0.FPCI_O\(69),
datad => \GRLFPC2_0.FPCI_O\(63),
datac => \GRLFPC2_0.FPCI_O\(70));
GRLFPC2_0_COMB_V_I_RDD_1_I_A3_15_5_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000f000f000f0")
port map (
combout => \GRLFPC2_0.COMB.V.I.RDD_1_I_A3_15_5_0\,
dataf => \GRLFPC2_0.FPCI_O\(47),
datae => \GRLFPC2_0.FPCI_O\(46),
datad => \GRLFPC2_0.FPCI_O\(45),
datac => \GRLFPC2_0.FPCI_O\(44));
GRLFPC2_0_COMB_V_I_RDD_1_I_A3_15_8: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000300000000")
port map (
combout => \GRLFPC2_0.COMB.V.I.RDD_1_I_A3_15_8\,
dataf => \GRLFPC2_0.COMB.V.I.RDD_1_I_A3_15_5_0\,
datae => \GRLFPC2_0.FPCI_O\(49),
datad => \GRLFPC2_0.FPCI_O\(48),
datac => \GRLFPC2_0.FPCI_O\(52),
datab => \GRLFPC2_0.FPCI_O\(50));
GRLFPC2_0_COMB_V_I_RDD_1_I_A3_15_7: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000ff")
port map (
combout => \GRLFPC2_0.COMB.V.I.RDD_1_I_A3_15_7\,
dataf => \GRLFPC2_0.FPCI_O\(59),
datae => \GRLFPC2_0.FPCI_O\(61),
datad => \GRLFPC2_0.FPCI_O\(51));
GRLFPC2_0_COMB_RDD_2_I_M3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff3000cfff0000")
port map (
combout => \GRLFPC2_0.N_83\,
dataf => \GRLFPC2_0.R.X.RDD\,
datae => \GRLFPC2_0.R.I.RDD\,
datad => N_37343_I_0,
datac => \GRLFPC2_0.R.I.V\,
datab => \GRLFPC2_0.R.I.EXEC\);
\GRLFPC2_0_COMB_V_I_PC_1_I_M2_23_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.N_3429\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.FPCI_O\(306),
datad => \GRLFPC2_0.R.I.PC_O\(23));
\GRLFPC2_0_WRADDR_1_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRADDRZ(1),
dataf => N_403,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.WRADDR_1_SQMUXA\,
datac => \GRLFPC2_0.R.I.INST\(27),
datab => N_356);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0ff00cccc")
port map (
combout => \GRLFPC2_0.N_3093\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => CPO_CCZ(0),
datac => N_676,
datab => N_612);
\GRLFPC2_0_COMB_DBGDATA_4_23_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(23),
dataf => \GRLFPC2_0.R.FSR.TEM\(0),
datae => N_400,
datad => N_401,
datac => N_689,
datab => N_625);
\GRLFPC2_0_COMB_V_I_PC_1_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.R.I.PC\(10),
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.FPCI_O\(293),
datad => \GRLFPC2_0.R.I.PC_O\(10));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcc3300fcfc3030")
port map (
combout => \GRLFPC2_0.N_3077\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.R.I.INST\(27),
datad => \GRLFPC2_0.FPCI_O\(310),
datac => \GRLFPC2_0.R.I.PC_O\(27),
datab => \GRLFPC2_0.N_91\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_70_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff000f0ffcc00cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(70),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.N_71\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_676,
datab => N_612);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_73_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0fff000ccffcc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(73),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.FPI.OP1\(39),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_676,
datab => N_612);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_257_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10503\,
dataf => \GRLFPC2_0.FPO.EXP\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_41_257_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff000f0ffcc00cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\(257),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.FPI.OP1\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_686,
datab => N_622);
GRLFPC2_0_COMB_UN1_V_STATE_RNIKKMB1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f30000000000")
port map (
combout => \GRLFPC2_0.N_1439\,
dataf => N_37318_1,
datae => \GRLFPC2_0.N_1015\,
datad => \GRLFPC2_0.COMB.V.STATE12_0\,
datac => \GRLFPC2_0.COMB.ISFPOP2_1\,
datab => \GRLFPC2_0.R.X.LD\);
GRLFPC2_0_COMB_UN1_FPCI_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => \GRLFPC2_0.N_1683\,
dataf => N_226,
datae => N_225);
GRLFPC2_0_COMB_UN3_HOLDN: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => \GRLFPC2_0.N_1685\,
dataf => N_157,
datae => N_156);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRONEMORE: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN12_SRTOSTICKY_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN12_SRTOSTICKY_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8_I\(57),
datad => N_53924,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3fcf00f030c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8_I\(57),
datae => N_53924,
datad => N_53884,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffff0000f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8_I\(57),
datae => N_53884,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3fcf00f030c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(32),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(31),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcf3f00f0c0300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(34),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(33),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_20_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff00f00cccccccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9994\,
dataf => \GRLFPC2_0.FPI.LDOP_0_1\,
datae => \GRLFPC2_0.FPI.OP2\(37),
datad => \GRLFPC2_0.FPI.OP2\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(136));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_20_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0cff0c00fcfffc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10114\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(20),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9994\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_37_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53946,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_20_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3fcf00f030c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(20),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(22),
datae => N_53946,
datad => N_53945,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_20_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ff333cc0cc000")
port map (
combout => N_54001,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(20),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(21),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_20_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00fff00f0fffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(20),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(20),
datae => N_54001,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff33fc30cf03cc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(27),
dataf => N_53879,
datae => N_53878,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(29),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(29),
datae => N_53879,
datad => N_53878,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(28),
dataf => N_53898,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3fcf0ff030c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(31),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(31),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(30),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(28),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53898,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ffffccf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(24),
dataf => N_53898,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ff333cc0cc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(24),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(24),
datae => N_53908,
datad => N_53903,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3fcc0cf333c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(25),
dataf => N_53879,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(25),
datad => N_53931,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_35_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffccf00000ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(35),
dataf => N_53877,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53886,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_40_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcffccc33033000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(40),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(38),
datae => N_53886,
datad => N_53885,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ffffccf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(29),
dataf => N_53896,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffccfcc33300300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(31),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(29),
datae => N_53878,
datad => N_53877,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_9_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcf3f00f0c0300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(9),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff0000f0f0f0f0")
port map (
combout => N_53938,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffc00fcff300030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(1),
dataf => N_53935,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datac => N_53938,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53984,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ffcc00f000cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(6),
dataf => N_53984,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53980,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53982,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcf3f00f0c0300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(6),
datae => N_53980,
datad => N_53982,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_21_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53885,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53919,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53890,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53889,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53887,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccfffff0cc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(32),
dataf => N_53887,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_30_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53878,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53877,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53896,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(33),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(33),
datae => N_53878,
datad => N_53877,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3fcf0ff030c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(33),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(33),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53945,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccfff0ffcc00f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(24),
dataf => N_53945,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53977,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_22_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffccfff000cc00f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(22),
dataf => N_53977,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_22_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(22),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(22),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(24),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53958,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53979,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_21_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcffccc33033000")
port map (
combout => N_54000,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(22),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(21),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_I\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_21_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cfc00f00fff03f30")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9817\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(36),
datae => N_54000,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIKDT6Q51_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(38),
dataf => N_27258,
datae => N_27278,
datad => N_27277);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIGTT7TL1_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(39),
dataf => N_27258,
datae => N_27280,
datad => N_27279);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fbf8cbc83b380b08")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10056\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(18),
datae => \GRLFPC2_0.FPO.FRAC\(38),
datad => \GRLFPC2_0.FPO.FRAC\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf3f0ff0c03000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(10),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(10),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(11),
dataf => N_53926,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffccfcc33300300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(13),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(11),
datae => N_53929,
datad => N_53874,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_15_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffccf3c03f0c3300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(15),
dataf => N_53929,
datae => N_53874,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffc3330cfcc0300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(17),
dataf => N_53874,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(15),
datad => N_53930,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_22_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcf3f0ff0c03000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(22),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(22),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_35_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53908,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_22_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcffccc33033000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(22),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(20),
datae => N_53908,
datad => N_53903,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53879,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_23_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffcffccc33033000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(23),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(21),
datae => N_53879,
datad => N_53931,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53904,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff3ff333cc0cc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(39),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(39),
datae => N_53892,
datad => N_53904,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffff0000f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8_I\(57),
datae => N_53905,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3fcf00f030c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8_I\(57),
datae => N_53875,
datad => N_53905,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8_I\(57),
datad => N_53875,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccff00f0f0f0f0")
port map (
combout => N_53884,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ccf0ffff0000")
port map (
combout => N_53905,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffccfcc33300300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(8),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(6),
datae => N_53875,
datad => N_53927,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ccf0ffff0000")
port map (
combout => N_53924,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(237));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccf0f0ff00ff00")
port map (
combout => N_53926,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(241));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccff00f0f0f0f0")
port map (
combout => N_53883,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(239));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ccf0ffff0000")
port map (
combout => N_53929,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(10),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(10),
datae => N_53875,
datad => N_53927,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccff00f0f0f0f0")
port map (
combout => N_53925,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(240));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(10),
dataf => N_53925,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffccfcc33300300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(12),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(10),
datae => N_53927,
datad => N_53907,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccff00f0f0f0f0")
port map (
combout => N_53927,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_14_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(14),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(14),
datae => N_53927,
datad => N_53907,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ffff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_14_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0ccfffff0cc0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(14),
dataf => N_53923,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_16_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffccfcc33300300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(16),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(14),
datae => N_53907,
datad => N_53895,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53880,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccf0ffffccf00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(39),
dataf => N_53880,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_20_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53892,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_16_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53891,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_41_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffccfcc33300300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(41),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(39),
datae => N_53892,
datad => N_53891,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_45_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53907,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(18),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(18),
datae => N_53907,
datad => N_53895,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_20_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff3ccc03f330c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(20),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(19),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(20),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRONEMORE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_43_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53923,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53903,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_41_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53895,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_20_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffccf00000ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(20),
dataf => N_53895,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_21_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcf3f00f0c0300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6_I\(21),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(20),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_40_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53930,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53931,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff33f33ccc00c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(19),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_I\(19),
datae => N_53874,
datad => N_53930,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1));
\GRLFPC2_0_COMB_RS2_1_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000fffff0000000")
port map (
combout => \GRLFPC2_0.COMB.RS2_1\(2),
dataf => \GRLFPC2_0.R.A.RS2\(2),
datae => N_13,
datad => \GRLFPC2_0.N_951\,
datac => N_55);
\GRLFPC2_0_COMB_DBGDATA_4_16_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => CPO_DBG_DATAZ(16),
dataf => \GRLFPC2_0.R.FSR.FTT\(2),
datae => N_400,
datad => N_401,
datac => N_682,
datab => N_618);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_16_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0ff00cccc")
port map (
combout => \GRLFPC2_0.N_3099\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.FSR.FTT\(2),
datac => N_682,
datab => N_618);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_14_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0ff00cccc")
port map (
combout => \GRLFPC2_0.N_3097\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.FSR.FTT\(0),
datac => N_680,
datab => N_616);
\GRLFPC2_0_WRADDR_1_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc0000f0cc")
port map (
combout => RFI2_WRADDRZ(3),
dataf => N_405,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => \GRLFPC2_0.WRADDR_1_SQMUXA\,
datac => \GRLFPC2_0.R.I.INST\(29),
datab => N_358);
\GRLFPC2_0_COMB_V_I_PC_1_I_M2_16_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.N_3423\,
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.FPCI_O\(299),
datad => \GRLFPC2_0.R.I.PC_O\(16));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00f0f0ff00cccc")
port map (
combout => \GRLFPC2_0.N_3091\,
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.R.A.AFSR\,
datad => \GRLFPC2_0.R.FSR.AEXC\(3),
datac => N_674,
datab => N_610);
GRLFPC2_0_COMB_WREN1_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000fc00fffffc00")
port map (
combout => RFI1_WRENZ,
dataf => N_401,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => N_13,
datac => \GRLFPC2_0.COMB.WREN1_9_IV_1\,
datab => \GRLFPC2_0.COMB.WREN1_9_IV_0\);
GRLFPC2_0_COMB_WREN2_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffc000000fc00")
port map (
combout => RFI2_WRENZ,
dataf => N_401,
datae => \GRLFPC2_0.WRADDR_0_SQMUXA_1\,
datad => N_13,
datac => \GRLFPC2_0.COMB.WREN2_9_IV_1\,
datab => \GRLFPC2_0.COMB.WREN2_9_IV_0\);
\GRLFPC2_0_COMB_V_I_PC_1_14_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.R.I.PC\(14),
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.FPCI_O\(297),
datad => \GRLFPC2_0.R.I.PC_O\(14));
\GRLFPC2_0_COMB_V_I_PC_1_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.R.I.PC\(8),
dataf => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
datae => \GRLFPC2_0.FPCI_O\(291),
datad => \GRLFPC2_0.R.I.PC_O\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_67_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0fff000ccffcc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(67),
dataf => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
datae => \GRLFPC2_0.N_71\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => N_682,
datab => N_618);
GRLFPC2_0_V_FSR_FTT_1_SQMUXA_I: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffccfffcff00fff0")
port map (
combout => \GRLFPC2_0.N_58\,
dataf => \GRLFPC2_0.N_76_I\,
datae => \GRLFPC2_0.R.X.LD\,
datad => \GRLFPC2_0.R.X.SEQERR\,
datac => \GRLFPC2_0.R.X.AFSR\,
datab => \GRLFPC2_0.R.X.AFQ\);
GRLFPC2_0_COMB_WREN2_9_IV_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffc00fc00fc00")
port map (
combout => \GRLFPC2_0.COMB.WREN2_9_IV_1\,
dataf => \GRLFPC2_0.WREN2_2_SQMUXA\,
datae => N_354,
datad => \GRLFPC2_0.WREN2_1_SQMUXA_0\,
datac => N_362,
datab => N_361);
GRLFPC2_0_COMB_WREN2_9_IV_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0cc00000000")
port map (
combout => \GRLFPC2_0.COMB.WREN2_9_IV_0\,
dataf => \GRLFPC2_0.N_1391\,
datae => \GRLFPC2_0.N_83\,
datad => \GRLFPC2_0.WRADDR_1_SQMUXA\,
datac => \GRLFPC2_0.R.I.INST\(25),
datab => N_354);
GRLFPC2_0_WREN2_1_SQMUXA_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000003000000000")
port map (
combout => \GRLFPC2_0.WREN2_1_SQMUXA_0\,
dataf => N_349,
datae => \GRLFPC2_0.R.X.SEQERR\,
datad => \GRLFPC2_0.N_1105\,
datac => \GRLFPC2_0.R.X.LD\,
datab => \GRLFPC2_0.R.X.AFSR\);
GRLFPC2_0_WREN2_2_SQMUXA: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000030")
port map (
combout => \GRLFPC2_0.WREN2_2_SQMUXA\,
dataf => \GRLFPC2_0.N_1105\,
datae => N_349,
datad => \GRLFPC2_0.R.X.SEQERR\,
datac => \GRLFPC2_0.R.X.LD\,
datab => \GRLFPC2_0.R.X.AFSR\);
GRLFPC2_0_COMB_WREN1_9_IV_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0300ffff03000300")
port map (
combout => \GRLFPC2_0.COMB.WREN1_9_IV_1\,
dataf => \GRLFPC2_0.WREN2_2_SQMUXA\,
datae => N_354,
datad => \GRLFPC2_0.WREN2_1_SQMUXA_0\,
datac => N_362,
datab => N_361);
GRLFPC2_0_COMB_ISFPOP2_1_0_M3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0ccf0f0f0f0f0")
port map (
combout => \GRLFPC2_0.COMB.ISFPOP2_1\,
dataf => \GRLFPC2_0.R.X.FPOP\,
datae => \GRLFPC2_0.R.I.EXEC\,
datad => \GRLFPC2_0.R.I.V\,
datac => \GRLFPC2_0.R.I.INST\(19),
datab => N_348);
GRLFPC2_0_R_I_V_RNIKA7K: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f030f030c000f000")
port map (
combout => \GRLFPC2_0.COMB.V.STATE12_0\,
dataf => \GRLFPC2_0.R.X.FPOP\,
datae => \GRLFPC2_0.R.X.SEQERR\,
datad => \GRLFPC2_0.R.I.EXEC\,
datac => \GRLFPC2_0.R.I.V\,
datab => \GRLFPC2_0.N_1105\);
\GRLFPC2_0_R_STATE_RNO_0_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000300000")
port map (
combout => \GRLFPC2_0.V.STATE_1_SQMUXA_3\,
dataf => \GRLFPC2_0.N_1015\,
datae => \GRLFPC2_0.N_76_I\,
datad => \GRLFPC2_0.R.X.SEQERR\,
datac => \GRLFPC2_0.R.X.AFQ\,
datab => \GRLFPC2_0.N_1105\);
GRLFPC2_0_COMB_QNE2_I_O3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.N_76_I\,
dataf => \GRLFPC2_0.R.STATE\(0),
datae => \GRLFPC2_0.R.STATE\(1));
GRLFPC2_0_COMB_UN1_FPCI_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff00")
port map (
combout => \GRLFPC2_0.N_1105\,
dataf => N_14,
datae => N_363,
datad => N_364);
GRLFPC2_0_COMB_WREN125: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000003000000000")
port map (
combout => \GRLFPC2_0.N_1391\,
dataf => N_37318_1,
datae => \GRLFPC2_0.R.X.LD\,
datad => \GRLFPC2_0.COMB.ISFPOP2_1\,
datac => \GRLFPC2_0.COMB.V.STATE12_0\,
datab => \GRLFPC2_0.N_1015\);
GRLFPC2_0_COMB_WREN1_9_IV_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0f3300000000")
port map (
combout => \GRLFPC2_0.COMB.WREN1_9_IV_0\,
dataf => \GRLFPC2_0.N_1391\,
datae => \GRLFPC2_0.N_83\,
datad => \GRLFPC2_0.WRADDR_1_SQMUXA\,
datac => \GRLFPC2_0.R.I.INST\(25),
datab => N_354);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TEMP\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0f000fff0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_64_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaaff00f0f0cccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(64),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
datad => \GRLFPC2_0.FPO.FRAC\(49),
datac => \GRLFPC2_0.FPO.FRAC\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => N_53935,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccff00f0f0f0f0")
port map (
combout => N_53875,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(238));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffafcfaff0a0c0a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10936\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN13_RESVEC\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(241));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000101ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10936\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10931\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7352\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM6\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_44_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => N_53874,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIQ83D_43_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10931\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_NORMDETECT_NOTSLFROMNORM_19_0_A2_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0c0f0f0c0f0c0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM12\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_X2_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => N_32762_I,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffc3000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_659\,
dataf => N_34180,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1714\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1736\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_1_A2_0_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1_A2_0\(39),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_1_O2_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffc000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8537\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1588\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1133\,
datad => N_32738_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1714\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1_A2_0\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O8_3_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f00300c00000c000")
port map (
combout => N_28243,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_PCTRL_1_CO5: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_4_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f000f0000000")
port map (
combout => N_28267,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O17_4_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff0000ffff000000")
port map (
combout => N_33061,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O17_4_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f000000f0f00f")
port map (
combout => N_33277,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O17_5_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000030c3000f000")
port map (
combout => N_33278,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_33368_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_X2_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => N_33547_I,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_X2_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => N_28892_I,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O23_7_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c000000030000f0")
port map (
combout => N_33565,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O9_2_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0f0f0fff000000")
port map (
combout => N_33769,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_X2_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => N_33798_I,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O22_5_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f000f00000000f")
port map (
combout => N_33813,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A2_12_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000000000")
port map (
combout => N_34007,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_X2_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => N_32959_I,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O23_2_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => N_34024,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_X2_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => N_34311_I,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O26_9_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff0000ffff00")
port map (
combout => N_34107,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_X2_0_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => N_34239_I,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_24_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_33721_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A11_0_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"03cc33ff00000000")
port map (
combout => N_28206,
dataf => N_33838_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_33734_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A14_5_2_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_32722_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_9_1_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_28652_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_11_1_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_32980_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_4_1_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_32908_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_5_1_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_34254_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A24_27_1_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_33144_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A23_1_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ff000000000000")
port map (
combout => N_33498_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_18_2_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000ff0000")
port map (
combout => N_33501_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_19_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000030000000000")
port map (
combout => N_33590,
dataf => N_33984_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_44_1_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_28250_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A3_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_33503_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A9_1_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3f000f0000000000")
port map (
combout => N_33778,
dataf => N_33735_1,
datae => N_33340_I,
datad => N_28222_1,
datac => N_33111,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O17_2_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => N_33055,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_X2_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => N_28681_I,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_1_1_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_29071_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_7_1_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_28251_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_33659_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_2_1_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_28212_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_9_1_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_28211_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_28_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_32786_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A26_22_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c00000000000000")
port map (
combout => N_33987,
dataf => N_28271_1,
datae => N_28564_2,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A22_1_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_28560_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_6_1_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_28227_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_10_1_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_32791_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_16_1_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_28549_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_O2_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_719\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_9_1_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_33447_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A32_10_1_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_28730_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_32723_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_19_1_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_28250_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A24_1_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_32731_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_0_1_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_33899_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A21_1_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_28492_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_9_1_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_28921_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_18_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_33543,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_16_1_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_34341_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_6_1_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_28658_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_O21_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_531\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A14_9_2_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_33140_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_5_1_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_32727_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_18_1_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_33574_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A14_4_1_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_32979_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A15_1_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_33146_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_3_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_29195_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A8_1_0_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_33577_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A19_1_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_33081_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_4_1_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_33138_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_7_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_33735_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_22_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_22__G2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8764\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9608\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9665\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9645\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9607\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_X2_1_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => N_33263_I,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_33074_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_8_2_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_32796_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_M27_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ffffffff00ff00")
port map (
combout => N_34233,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_M3_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0cf0f3ff00f0f")
port map (
combout => N_33411,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_14_2_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_33507_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_O28_0_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ffffffff")
port map (
combout => N_33178,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_O23_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffffffff")
port map (
combout => N_33548,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_2_1_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_28222_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_1_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_29366_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_3_1_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_28261_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A11_4_1_61_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_32844_3,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_3_1_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_32982_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_6_1_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_29518_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A14_5_1_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_28634_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_32844_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O2_0_0_O2_62_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000c00000300033")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8524\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_0_O2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0fffffff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_479\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(71),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(74),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNILFOV1_248_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffff0fcf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_893\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_I_O2_3_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_O2_2_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00030000ffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1846\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_429\,
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_55_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f0fff000f000f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5330\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(12),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(60));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI85KHTB_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_176__G2\,
dataf => N_27258,
datae => N_27312,
datad => N_27311);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIC1OBQG_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(54),
dataf => N_27258,
datae => N_27310,
datad => N_27309);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIKUAVFK1_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(52),
dataf => N_27258,
datae => N_27306,
datad => N_27305);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIGVPO8J2_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(53),
dataf => N_27258,
datae => N_27308,
datad => N_27307);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI4Q19IP2_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(49),
dataf => N_27258,
datae => N_27300,
datad => N_27299);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI8EJI351_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(51),
dataf => N_27258,
datae => N_27304,
datad => N_27303);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIKOLUL62_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(47),
dataf => N_27258,
datae => N_27296,
datad => N_27295);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI4M7CDT_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(50),
dataf => N_27258,
datae => N_27302,
datad => N_27301);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNIO3FNKN3_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.FPO.FRAC\(48),
dataf => N_27258,
datae => N_27298,
datad => N_27297);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CHECKOVANDDENORM_UN13_NOTPOSSIBLEOV: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"8000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\,
dataf => \GRLFPC2_0.FPO.FRAC\(54),
datae => \GRLFPC2_0.FPO.FRAC\(52),
datad => \GRLFPC2_0.FPO.FRAC\(53),
datac => \GRLFPC2_0.FPO.FRAC\(49),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_16_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000fffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1503\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_547\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_O2_11_RNIBGS11_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1839\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_492\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1618\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNICKCS1_233_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffcffff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1544\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1839\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_429\,
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_O2_10_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_446\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_2_I_O2_10_4\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(255),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(254),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(256));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIEP39_247_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_I_O2_3_0\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(247),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(249));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_O2_17_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_547\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_A2_28_RNIRB3G2_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0300ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1852\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_893\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_389\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1636\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_I_O2_3_0\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIAU7Q_46_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00f000f000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1618\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_12_RNIN8TC5_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffcccc00c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1544\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1852\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1503\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1633\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1618\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_27_D_S_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ff0000000000")
port map (
combout => N_44786,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(51),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(50),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI0TSKGE3_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2\,
dataf => N_27316,
datae => N_27258,
datad => N_27315);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNI4DCT32_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_175__G2\,
dataf => N_27258,
datae => N_27314,
datad => N_27313);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_25_D: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0c3c3c3f0f0c3f0")
port map (
combout => N_44753,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(51));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_14: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ddd788827d772822")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10909\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10905\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.CONDITIONAL\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(51));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_7: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c999c39369396333")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10902\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(12),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SFTLFT.AREGXORBREG\,
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(51));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_27_D_D_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fdb97531eca86420")
port map (
combout => N_44787,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10902\,
datae => N_44753,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10911\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10909\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(50));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_27_D_D_0_RNIQUBP2R2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000200010003")
port map (
combout => D_N_7,
dataf => N_44787,
datae => N_53932,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_663\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK\,
dataa => N_44786);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTABORTNULLEXC: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ff00ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN25_LOCOV_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.REEXCOVUV.UN25_LOCOV_0\,
dataf => \GRLFPC2_0.FPO.EXP\(9),
datae => \GRLFPC2_0.FPO.EXP\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_24_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cc00cc000c000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1566\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_426\,
datae => N_33718_1,
datad => N_32738_1_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(67));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_2_1_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_34329_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_5_1_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_32782_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_257_RNI2N0G5: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_33725_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_1_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_33607_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_5_0_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_33652_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_12_1_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_28264_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN13_LOCOV_4: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.REEXCOVUV.UN13_LOCOV_4\,
dataf => \GRLFPC2_0.FPO.EXP\(6),
datae => \GRLFPC2_0.FPO.EXP\(5),
datad => \GRLFPC2_0.FPO.EXP\(4),
datac => \GRLFPC2_0.FPO.EXP\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN13_LOCOV_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.REEXCOVUV.UN13_LOCOV_3\,
dataf => \GRLFPC2_0.FPO.EXP\(7),
datae => \GRLFPC2_0.FPO.EXP\(2),
datad => \GRLFPC2_0.FPO.EXP\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN18_LOCOV: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5335\,
dataf => \GRLFPC2_0.FPO.EXP\(10),
datae => \GRLFPC2_0.FPO.EXP\(9),
datad => \GRLFPC2_0.FPO.EXP\(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_16_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00000000ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10911\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_10: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f00ff0f00f0f0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10905\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_AREGXORBREG_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SFTLFT.AREGXORBREG\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_CONDITIONAL_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.CONDITIONAL\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_O2_12_4_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_O2_12_4\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(238),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(241),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(240),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(239));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_O2_12_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_504\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_O2_12_4\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(237));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNID7UL_234_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffcffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_I_O2_0\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_O2_11_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff3fffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_492\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_O2_11_3\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(238),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(241),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(239),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(240));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIJ9LD_234_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ffffffffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_429\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_O2_11_RNIC8VE1_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffc0ffcc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_770\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_492\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_429\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_I_O2_0\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_12_RNI07NV1_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff00030000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_770\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1633\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_49_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(49),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_40_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(40),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_39_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(39),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_30_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ff0000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(30),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_44_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(44),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_32_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(32),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_54_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(54),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(36),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_50: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"1428000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_50\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_42\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_28\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(49),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(40));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_52_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(52),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_35_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(35),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(53),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_34_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(34),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_27_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ff0000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(27),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_26_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ff0000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(26),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ff0000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(25),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ff0000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(10),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_16: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f00f00f00f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_16\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(10),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(25));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(56),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_37_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(37),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_46_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(46),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0000000f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(31),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_47_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(47),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_38_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(38),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(51),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_43_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(43),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_20_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ff0000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(20),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ff0000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(13),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_7: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f00f00f00f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(13),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(20),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(20));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_24_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0ff00f0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(24),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_21_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ff0000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(21),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_6: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f00f00f00f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(21),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(24),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffc000000fc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(115),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN38_SHDVAR_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5416\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffc000000fc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000033003300000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5391\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5410\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_29_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ff0000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(29),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_45_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(45),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(57),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f00ff00fcc3300ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(57),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(174));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_28_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ff0000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(28),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0ff00f0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_15_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ff0000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(15),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0ff00f0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_14: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f00f00f00f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_14\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(15),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_23_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ff0000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(23),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_14_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0ff00f0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(14),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_22_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0ff00f0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(22),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_12: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f00f00f00f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_12\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(22),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_18_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ff0000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(18),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ff0000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(11),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ff0000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(19),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0ff00f0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(8),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_10: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f00f00f00f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_10\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(19),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ff0000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(17),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_9_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0ff00f0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(9),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_16_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ff0000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(16),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0ff0000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_8: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f00f00f00f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(16),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(16));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_33: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"030c30c000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_33\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_8\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_46: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"1248000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_46\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_33\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_10\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(48),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(42),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_50_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(50),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_41_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(41),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_55_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff000000ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(55),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(33),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0ff00f0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffc000000fc00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0ff00f0f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(12),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_5: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0110022004400880")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(12),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_51: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"1248000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_51\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_44\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_XZXBUS\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(33));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"8000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_53\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_51\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_50\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_46\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_48\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_47\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10871\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(256));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10870\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(257));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_9_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33ccff000ff0ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(9),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_9_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10879\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33ccff000ff0ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(8),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10878\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(249));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff03cf0f0f03cf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(238));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10876\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(238),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(251));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff03cf0f0f03cf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(6),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(239));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10875\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(239),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(252));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5339\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(232));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_12_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10882\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(232),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(245));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5301\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10880\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(247));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5343\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10881\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff0ff0033ccff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(240));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10874\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(240),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(253));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_1_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10861\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33ccff000ff0ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(237),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10877\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(250),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(237));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_5: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffffeb")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_7\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10873\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(241),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(254));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_COMPUTECONST_UN13_RESVEC: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN13_RESVEC\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_8: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffd8ff27")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_6\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10860\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10873\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10872\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(255));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_NE: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffd8ff27")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_10\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10859\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10872\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_333_RNIVPQS3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_34263_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A14_1_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_28857_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_33070_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A26_12_0_11_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A26_12_0\(11),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_30_1_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_28564_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_X2_48_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => N_33340_I,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_32_RNIQ9HN5: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11641\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O23_3_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffffffff")
port map (
combout => N_34029,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_10_0_A2_RNII7KE1_60_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c000c000cc00c000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1568\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_603\,
datae => N_34029,
datad => N_33340_I,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9509\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_11_0_O2_RNIK29P9_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0f0fffff0003")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_458\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3945_I_I_O2_3_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1568\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_473\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_25_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1730\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_458\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(67));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A9_1_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_29262_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_2_1_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_28266_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_7_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_32738_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_13_1_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_28271_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A23_1_31_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_32730_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_5_1_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_32909_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_4_2_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_33297_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_O2_53_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_797\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_32738_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O25_11_19_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_782\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_0_0_O2_56_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000ffff")
port map (
combout => N_33179,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O32_9_57_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffffffff")
port map (
combout => N_33111,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O15_0_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => N_33004,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_33984_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_333_RNIC4NC1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_604\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_X2_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffff0000")
port map (
combout => N_32818_I,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O14_6_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00ffff00ff00ffff")
port map (
combout => N_53933,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_12_2_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_33436_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_4_2_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => N_29653_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O14_1_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffffffff")
port map (
combout => N_32821,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_51_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_32861_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O20_0_36_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_603\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_4_1_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffff00000000")
port map (
combout => N_32859_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A23_1_59_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => N_32858_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O14_4_25_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f00000ff000f000")
port map (
combout => N_32831,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_0_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_410\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_O24_33_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000ffffffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_419\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_1_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_RESULT_IV_0_RNI5I481_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0fffff030fffff")
port map (
combout => N_65584,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE\(12),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_0\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_20_RNIV70L: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f00000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
dataf => \GRLFPC2_0.FPI.LDOP_I_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_RETO\,
datad => RFO2_DATA1_RETO(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(95));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_19_RNIA80L: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f00000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
dataf => \GRLFPC2_0.FPI.LDOP_I_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_RETO\,
datad => RFO2_DATA1_RETO(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(94));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_18_RNI780L: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f00000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
dataf => \GRLFPC2_0.FPI.LDOP_I_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_RETO\,
datad => RFO2_DATA1_RETO(20),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(92));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_5_RNIUADH: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f00000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
dataf => \GRLFPC2_0.FPI.LDOP_I_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_RETO\,
datad => RFO2_DATA1_RETO(22),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(90));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_21_RNIT70L: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f00000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
dataf => \GRLFPC2_0.FPI.LDOP_I_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_RETO\,
datad => RFO2_DATA1_RETO(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(96));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_16_RNI380L: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f00000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
dataf => \GRLFPC2_0.FPI.LDOP_I_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_RETO\,
datad => RFO2_DATA1_RETO(24),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(88));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_15_RNI480L: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f00000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
dataf => \GRLFPC2_0.FPI.LDOP_I_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_RETO\,
datad => RFO2_DATA1_RETO(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(89));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_17_RNI880L: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f00000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
dataf => \GRLFPC2_0.FPI.LDOP_I_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_RETO\,
datad => RFO2_DATA1_RETO(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(87));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_23_RNI280L: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f00000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
dataf => \GRLFPC2_0.FPI.LDOP_I_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_RETO\,
datad => RFO2_DATA1_RETO(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(97));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_24_RNI180L: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f00000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
dataf => \GRLFPC2_0.FPI.LDOP_I_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_RETO\,
datad => RFO2_DATA1_RETO(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(98));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_25_RNI580L: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f00000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
dataf => \GRLFPC2_0.FPI.LDOP_I_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_RETO\,
datad => RFO2_DATA1_RETO(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(99));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_26_RNI880L: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f00000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
dataf => \GRLFPC2_0.FPI.LDOP_I_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_RETO\,
datad => RFO2_DATA1_RETO(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(100));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_27_RNIB80L: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f00000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102),
dataf => \GRLFPC2_0.FPI.LDOP_I_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_RETO\,
datad => RFO2_DATA1_RETO(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(102));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_60_RNI580L: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f00000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
dataf => \GRLFPC2_0.FPI.LDOP_I_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_RETO\,
datad => RFO2_DATA1_RETO(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(104));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_62_RNI880L: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f00000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
dataf => \GRLFPC2_0.FPI.LDOP_I_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_RETO\,
datad => RFO2_DATA1_RETO(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(105));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_30_RNI280L: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f00000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
dataf => \GRLFPC2_0.FPI.LDOP_I_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_RETO\,
datad => RFO2_DATA1_RETO(28),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(84));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_31_RNI080L: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f00000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
dataf => \GRLFPC2_0.FPI.LDOP_I_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_RETO\,
datad => RFO2_DATA1_RETO(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(86));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_33_RNI580L: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f00000ff000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
dataf => \GRLFPC2_0.FPI.LDOP_I_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_RETO\,
datad => RFO2_DATA1_RETO(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(85));
N_66969 <= not N_59;
N_66970 <= not \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42);
N_66971 <= not \GRLFPC2_0.FPI.LDOP_0_0\;
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
d => N_66446,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
d => N_66445,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4),
d => N_66444,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_91: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_141_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(141),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(141),
clk => N_12,
clrn => VCC,
ena => N_61580,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_13_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(13),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7248\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_248_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(248),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_246_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(246),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_249_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(249),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(249),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_247_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(247),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(247),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_29_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(29),
clk => N_12,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_30_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(30),
clk => N_12,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_233_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233),
d => N_37423,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_234_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234),
d => N_37230,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_236_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236),
d => N_37176,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_235_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235),
d => N_37203,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_251_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(251),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(251),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_253_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(253),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(253),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_257_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(257),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(257),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_252_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(252),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(252),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_80: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_I_O2_4_4\(4),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_I_O2_4_4_RETI\(4),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_250_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(250),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(250),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_255_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(255),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(255),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_254_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(254),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(254),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_130: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1_RETO\(115),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(115),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_111: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0_RETO\(71),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(71),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_110: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1_RETO\(71),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(71),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_45: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO\(3),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M\(3),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_3: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO\(1),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M\(1),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_37: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_90: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => N_65609_RETO,
d => N_65609,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_46: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_7: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_242_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242),
d => N_37417,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_243_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243),
d => N_37416,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_237_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(237),
d => N_37422,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_135: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(72),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(72),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_97: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(60),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(60),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_92: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(59),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(59),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_8: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_244_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244),
d => N_37415,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_256_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(256),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(256),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_241_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(241),
d => N_37418,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_240_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(240),
d => N_37419,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_239_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(239),
d => N_37420,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_238_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(238),
d => N_37421,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_232_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(232),
d => N_37424,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_245_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(245),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(245),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(4),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4424\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_7_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW\(7),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_43: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_BUSY_RET: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPO.BUSY_O\,
d => \GRLFPC2_0.R.MK.BUSY_RET_0_0_G0_MUX2\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_14: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_61_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(61),
clk => N_12,
clrn => VCC,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(61),
sload => N_66971,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_42: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5346\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5346_RETI\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(15),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_15__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_231_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(231),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(0),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_62_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(62),
clk => N_12,
clrn => VCC,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(62),
sload => N_66971,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_57_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10017\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10077\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_64: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(84),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(84),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_73: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(85),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(85),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_70: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(86),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(86),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_62: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(105),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(105),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_60: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(104),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(104),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_58: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(102),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(102),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_141: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(80),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(80),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_138: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(79),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(79),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_56: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(100),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(100),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_127: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(64),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(64),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_54: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(99),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(99),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_51: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(98),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(98),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_53: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(97),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(97),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_45: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(89),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(89),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_47: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(87),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(87),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_43: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(88),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(88),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_41: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(96),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(96),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_39: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(90),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(90),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_35: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(95),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(95),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_124: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(77),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(77),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_36: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(92),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(92),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_38: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(94),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(94),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_82_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(82),
clk => N_12,
clrn => VCC,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(82),
sload => N_66971,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_121: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(76),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(76),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_78_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(78),
clk => N_12,
clrn => VCC,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(78),
sload => N_66971,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_81_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(81),
clk => N_12,
clrn => VCC,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(81),
sload => N_66971,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_118: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(74),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(74),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_68_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(68),
clk => N_12,
clrn => VCC,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(68),
sload => N_66971,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_67_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(67),
clk => N_12,
clrn => VCC,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(67),
sload => N_66971,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_75_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(75),
clk => N_12,
clrn => VCC,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(75),
sload => N_66971,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_73_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(73),
clk => N_12,
clrn => VCC,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(73),
sload => N_66971,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_66_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(66),
clk => N_12,
clrn => VCC,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(66),
sload => N_66971,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_65_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(65),
clk => N_12,
clrn => VCC,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(65),
sload => N_66971,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_70_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(70),
clk => N_12,
clrn => VCC,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(70),
sload => N_66971,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_69_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(69),
clk => N_12,
clrn => VCC,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(69),
sload => N_66971,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_83_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(83),
clk => N_12,
clrn => VCC,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(83),
sload => N_66971,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_63_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(63),
clk => N_12,
clrn => VCC,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(63),
sload => N_66971,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_I\ <= not \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462\;
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_111_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(111),
clk => N_12,
clrn => VCC,
asdata => N_667,
sclr => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_I\,
sload => \GRLFPC2_0.FPI.LDOP\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_110_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(110),
clk => N_12,
clrn => VCC,
asdata => N_668,
sclr => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_I\,
sload => \GRLFPC2_0.FPI.LDOP\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_107_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(107),
clk => N_12,
clrn => VCC,
asdata => N_671,
sclr => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_I\,
sload => \GRLFPC2_0.FPI.LDOP\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_106_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(106),
clk => N_12,
clrn => VCC,
asdata => N_672,
sclr => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_I\,
sload => \GRLFPC2_0.FPI.LDOP\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_103_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(103),
clk => N_12,
clrn => VCC,
asdata => N_675,
sclr => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_I\,
sload => \GRLFPC2_0.FPI.LDOP\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_101_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(101),
clk => N_12,
clrn => VCC,
asdata => N_677,
sclr => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_I\,
sload => \GRLFPC2_0.FPI.LDOP\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_93_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(93),
clk => N_12,
clrn => VCC,
asdata => N_685,
sclr => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_I\,
sload => \GRLFPC2_0.FPI.LDOP\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_91_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(91),
clk => N_12,
clrn => VCC,
asdata => N_687,
sclr => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_I\,
sload => \GRLFPC2_0.FPI.LDOP\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_112_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(112),
clk => N_12,
clrn => VCC,
asdata => N_666,
sclr => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_I\,
sload => \GRLFPC2_0.FPI.LDOP\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_142: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(80),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(80),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_140: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPI.LDOP_RETO\,
d => \GRLFPC2_0.FPI.LDOP_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_139: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(79),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(79),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_137: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(72),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(72),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_136: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_132: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0_RETO\(115),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(115),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_128: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(64),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(64),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_125: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(77),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(77),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_122: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(76),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(76),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_119: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(74),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(74),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_116: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(72),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(72),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_114: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(71),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(71),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_112: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_108: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(71),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(71),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_97: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_96: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_95: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_94: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => D_N_7_RETO,
d => D_N_7,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => N_65488_RETO,
d => N_65488,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_2: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_105: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_372__G1_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_372__G1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_102: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(113),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(113),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_32_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_31_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_43_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(43),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_101: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPI.RST_1_RETO\,
d => \GRLFPC2_0.FPI.RST_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_100: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPI.LDOP_1_RETO\,
d => \GRLFPC2_0.FPI.LDOP_1_2\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_99: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_319__G1_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_319__G1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_BUSY_RET_1: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => RST_RETO,
d => N_11,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_44: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(9),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2_RETI\(9),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_RETI\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_36: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349_RETI\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_227_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(227),
d => \GRLFPC2_0.FPO.FRAC\(4),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_229_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(229),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(2),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_94: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_318__G1_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_318__G1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_90: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(51),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_89: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPO.FRAC_RETO\(4),
d => \GRLFPC2_0.FPO.FRAC\(4),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_11: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => N_59000_RETO,
d => N_59000,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_85: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_RETO\(50),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_84: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPO.FRAC_RETO\(5),
d => \GRLFPC2_0.FPO.FRAC\(5),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_83: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => N_58999_RETO,
d => N_58999,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_82: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_8: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => N_59001_RETO,
d => N_59001,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_79: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_3_I_RETO\(0),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_3_I\(0),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_78: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0_RETO\(114),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(114),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_76: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1_RETO\(114),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(114),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_92: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO(7),
d => N_60,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_86: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_85: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(55),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_30: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(80),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_78: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(53),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_24: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(78),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_74: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(54),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_70: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO5_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO5\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_68: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO(9),
d => N_62,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_67: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_65: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_TZ_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_TZ\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_0: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_58: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(85),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_57: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_55: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(0),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT\(0),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_53: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(56),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(56),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_52: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_49: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC_RETI\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_48: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO(11),
d => N_64,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7352\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7352_RETI\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_3__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_5_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_5__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_7_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_7__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_9_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_9__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_8_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_8__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_4: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM6\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM6_RETI\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_33: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => RFO2_DATA1_RETO(27),
d => N_693,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_31: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => RFO2_DATA1_RETO(26),
d => N_692,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_30: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => RFO2_DATA1_RETO(28),
d => N_694,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_29: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => RFO2_DATA1_RETO(7),
d => N_673,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_28: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => RFO2_DATA1_RETO(8),
d => N_674,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_27: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => RFO2_DATA1_RETO(10),
d => N_676,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_26: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => RFO2_DATA1_RETO(12),
d => N_678,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_25: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => RFO2_DATA1_RETO(13),
d => N_679,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_24: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => RFO2_DATA1_RETO(14),
d => N_680,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_23: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => RFO2_DATA1_RETO(15),
d => N_681,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_17: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => RFO2_DATA1_RETO(25),
d => N_691,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_49: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPI.LDOP_I_RETO\,
d => N_66971,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_15: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => RFO2_DATA1_RETO(23),
d => N_689,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_16: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => RFO2_DATA1_RETO(24),
d => N_690,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_21: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => RFO2_DATA1_RETO(16),
d => N_682,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_5: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => RFO2_DATA1_RETO(22),
d => N_688,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_18: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => RFO2_DATA1_RETO(20),
d => N_686,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_19: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => RFO2_DATA1_RETO(18),
d => N_684,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_12: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7350\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7350_RETI\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_13_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_13__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_12_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_12__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_11_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_11__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_14_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_14__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_9: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_0_RETI\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_16_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_16__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_6_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_6__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(11),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(11),
clk => N_12,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_374_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(374),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(374),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(9),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(9),
clk => N_12,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(12),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(12),
clk => N_12,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_15__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_17_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_17__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_34: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5\(2),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5_RETI\(2),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_20: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => RFO2_DATA1_RETO(17),
d => N_683,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_0: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_6: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => RFO2_DATA1_RETO(3),
d => N_669,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_1: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => RFO2_DATA1_RETO(4),
d => N_670,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_7: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_3\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_3_RETI\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_10__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_3: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => N_65775,
d => N_65775_RETI,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_2: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => N_65496,
d => N_65496_RETI,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_41: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_40: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_39: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_16_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(10),
clk => N_12,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(1),
clk => N_12,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_376_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(376),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_DIVMULTV\(0),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_14_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(14),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(14),
clk => N_12,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_35: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO(5),
d => N_58,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_34: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_29: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO(12),
d => N_65,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_28: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(84),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_23: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO(8),
d => N_61,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_22: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_17: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO(10),
d => N_63,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_16: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_15: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_11: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(81),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_10: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_5: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_4: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_375_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(375),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(375),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_13_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(13),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(13),
clk => N_12,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_I_V: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.V\,
d => N_38488,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_67_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(67),
d => N_38487,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_63_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(63),
d => \GRLFPC2_0.COMB.V.I.RES_1\(63),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_59_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(59),
d => \GRLFPC2_0.FPO.EXP\(7),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(62),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_58_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(58),
d => \GRLFPC2_0.FPO.EXP\(6),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(61),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_57_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(57),
d => \GRLFPC2_0.FPO.EXP\(5),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(60),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_56_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(56),
d => \GRLFPC2_0.FPO.EXP\(4),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(59),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_55_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(55),
d => \GRLFPC2_0.FPO.EXP\(3),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(58),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_54_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(54),
d => \GRLFPC2_0.FPO.EXP\(2),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(57),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_53_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(53),
d => \GRLFPC2_0.FPO.EXP\(1),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(56),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_52_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(52),
d => \GRLFPC2_0.FPO.EXP\(0),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(55),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_51_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(51),
d => \GRLFPC2_0.FPO.FRAC\(54),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(54),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_50_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(50),
d => \GRLFPC2_0.FPO.FRAC\(53),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(53),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_49_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(49),
d => \GRLFPC2_0.FPO.FRAC\(52),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(52),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_48_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(48),
d => \GRLFPC2_0.FPO.FRAC\(51),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(51),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_47_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(47),
d => \GRLFPC2_0.FPO.FRAC\(50),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(50),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_46_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(46),
d => \GRLFPC2_0.FPO.FRAC\(49),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(49),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_45_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(45),
d => \GRLFPC2_0.FPO.FRAC\(48),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(48),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_44_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(44),
d => \GRLFPC2_0.FPO.FRAC\(47),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(47),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_43_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(43),
d => \GRLFPC2_0.FPO.FRAC\(46),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(46),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_42_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(42),
d => \GRLFPC2_0.FPO.FRAC\(45),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(45),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_41_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(41),
d => \GRLFPC2_0.FPO.FRAC\(44),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(44),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_40_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(40),
d => \GRLFPC2_0.FPO.FRAC\(43),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(43),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_39_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(39),
d => \GRLFPC2_0.FPO.FRAC\(42),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(42),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_38_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(38),
d => \GRLFPC2_0.FPO.FRAC\(41),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(41),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_37_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(37),
d => \GRLFPC2_0.FPO.FRAC\(40),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(40),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_36_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(36),
d => \GRLFPC2_0.FPO.FRAC\(39),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(39),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_35_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(35),
d => \GRLFPC2_0.FPO.FRAC\(38),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(38),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_34_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(34),
d => \GRLFPC2_0.FPO.FRAC\(37),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(37),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_33_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(33),
d => \GRLFPC2_0.FPO.FRAC\(36),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(36),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_32_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(32),
d => \GRLFPC2_0.FPO.FRAC\(35),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(35),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_31_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(31),
d => \GRLFPC2_0.FPO.FRAC\(34),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(34),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_30_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(30),
d => \GRLFPC2_0.FPO.FRAC\(33),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(33),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_29_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(29),
d => \GRLFPC2_0.FPO.FRAC\(32),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
asdata => \GRLFPC2_0.FPI.OP2\(32),
sload => \GRLFPC2_0.N_1438\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_116_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(116),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2\,
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(118),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_117_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(117),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_175__G2\,
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(119),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_118_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(118),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_176__G2\,
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(120),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_119_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(119),
d => \GRLFPC2_0.FPO.FRAC\(54),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(121),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_120_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(120),
d => \GRLFPC2_0.FPO.FRAC\(53),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(122),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_121_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(121),
d => \GRLFPC2_0.FPO.FRAC\(52),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(123),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_122_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(122),
d => \GRLFPC2_0.FPO.FRAC\(51),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(124),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_123_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(123),
d => \GRLFPC2_0.FPO.FRAC\(50),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(125),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_124_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(124),
d => \GRLFPC2_0.FPO.FRAC\(49),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(126),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_125_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(125),
d => \GRLFPC2_0.FPO.FRAC\(48),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(127),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_126_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(126),
d => \GRLFPC2_0.FPO.FRAC\(47),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(128),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_127_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(127),
d => \GRLFPC2_0.FPO.FRAC\(46),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(129),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_128_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(128),
d => \GRLFPC2_0.FPO.FRAC\(45),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(130),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_129_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(129),
d => \GRLFPC2_0.FPO.FRAC\(44),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(131),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_130_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(130),
d => \GRLFPC2_0.FPO.FRAC\(43),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(132),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_131_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(131),
d => \GRLFPC2_0.FPO.FRAC\(42),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(133),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_132_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(132),
d => \GRLFPC2_0.FPO.FRAC\(41),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(134),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_133_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(133),
d => \GRLFPC2_0.FPO.FRAC\(40),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(135),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_134_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(134),
d => \GRLFPC2_0.FPO.FRAC\(39),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(136),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_135_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(135),
d => \GRLFPC2_0.FPO.FRAC\(38),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(137),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_136_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(136),
d => \GRLFPC2_0.FPO.FRAC\(37),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(138),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_137_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(137),
d => \GRLFPC2_0.FPO.FRAC\(36),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(139),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_138_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(138),
d => \GRLFPC2_0.FPO.FRAC\(35),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(140),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_139_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(139),
d => \GRLFPC2_0.FPO.FRAC\(34),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(141),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_140_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(140),
d => \GRLFPC2_0.FPO.FRAC\(33),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(142),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_142_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(142),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(142),
clk => N_12,
clrn => VCC,
ena => N_61580,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_143_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(143),
d => \GRLFPC2_0.FPO.FRAC\(30),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(145),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_144_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(144),
d => \GRLFPC2_0.FPO.FRAC\(29),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(146),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_145_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(145),
d => \GRLFPC2_0.FPO.FRAC\(28),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(147),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_146_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(146),
d => \GRLFPC2_0.FPO.FRAC\(27),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(148),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_147_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(147),
d => \GRLFPC2_0.FPO.FRAC\(26),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(149),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_148_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(148),
d => \GRLFPC2_0.FPO.FRAC\(25),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(150),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_149_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(149),
d => \GRLFPC2_0.FPO.FRAC\(24),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(151),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_150_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(150),
d => \GRLFPC2_0.FPO.FRAC\(23),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(152),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_151_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(151),
d => \GRLFPC2_0.FPO.FRAC\(22),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(153),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_152_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(152),
d => \GRLFPC2_0.FPO.FRAC\(21),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(154),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_153_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(153),
d => \GRLFPC2_0.FPO.FRAC\(20),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(155),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_154_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(154),
d => \GRLFPC2_0.FPO.FRAC\(19),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(156),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_155_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(155),
d => \GRLFPC2_0.FPO.FRAC\(18),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(157),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_156_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(156),
d => \GRLFPC2_0.FPO.FRAC\(17),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(158),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_157_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(157),
d => \GRLFPC2_0.FPO.FRAC\(16),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(159),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_158_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(158),
d => \GRLFPC2_0.FPO.FRAC\(15),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(160),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_159_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(159),
d => \GRLFPC2_0.FPO.FRAC\(14),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(161),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_160_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(160),
d => \GRLFPC2_0.FPO.FRAC\(13),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(162),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_161_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(161),
d => \GRLFPC2_0.FPO.FRAC\(12),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(163),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_162_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(162),
d => \GRLFPC2_0.FPO.FRAC\(11),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(164),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_163_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(163),
d => \GRLFPC2_0.FPO.FRAC\(10),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(165),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_164_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(164),
d => \GRLFPC2_0.FPO.FRAC\(9),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(166),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_165_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(165),
d => \GRLFPC2_0.FPO.FRAC\(8),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(167),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_166_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(166),
d => \GRLFPC2_0.FPO.FRAC\(7),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(168),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_167_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(167),
d => \GRLFPC2_0.FPO.FRAC\(6),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(169),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_168_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(168),
d => \GRLFPC2_0.FPO.FRAC\(5),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(170),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_169_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(169),
d => \GRLFPC2_0.FPO.FRAC\(4),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(171),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_170_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(170),
d => \GRLFPC2_0.FPO.FRAC\(3),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(172),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_171_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(171),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(2),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_14\(171),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_172_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(172),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(1),
clk => N_12,
clrn => VCC,
ena => N_61580,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_14\(172),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10373_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_77_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_49_I\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_76_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7272\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_74_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(74),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7274\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_73_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_51_I\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_72_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_71_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(71),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.UN36_PCTRL_NEW_I\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_70_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(70),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(68),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_68_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(68),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3926\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_66_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(66),
d => \GRLFPC2_0.FPI.START\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_65_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW_2\(65),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_64_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(64),
d => \GRLFPC2_0.FPI.RST\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_63_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(63),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_62_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(62),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_61_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(61),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__I0_I_2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_60_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(60),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_59_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(59),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_58_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(58),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_57_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(57),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_57__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_56_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(56),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_55_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(55),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_54_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(54),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_53_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(53),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_52_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_51_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(51),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_50_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(50),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_49_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(49),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_48_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_48__I0_I_0\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_47_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(47),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_47__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_46_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(46),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_46__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_45_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_44_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_44__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_42_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_41_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(41),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_41__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_40_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(40),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_40__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_39_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(39),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_39__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_38_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(38),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_16_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(16),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SCTRL_NEW\(0),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
d => N_66970,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_14_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(14),
d => N_53873,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_12_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_I_I_0\(0),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_11_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
d => N_66969,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_9_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(9),
d => N_36985,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_8_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(8),
d => N_36986,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_6_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(6),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4459\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_5_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(5),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4465_I\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(3),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4874\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(2),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7259\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(1),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7260\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(0),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW_6\(0),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_36_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_35_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(35),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_35__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_34_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_33_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_28_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_27_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_26_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_25_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_24_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(24),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_24__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_23_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(23),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_23__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_22_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(22),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_22__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_21_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(21),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_21__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_20_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(20),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_20__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_19_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(19),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_18_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(18),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(8),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_8__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(5),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(2),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_2__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(1),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_1__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_377_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(377),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF\(0),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_373_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(373),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_3_I\(0),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_372_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(372),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_372__G1\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_371_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(371),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(112),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_370_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(370),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(111),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_369_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(369),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(110),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_368_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(368),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(109),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_367_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(367),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(108),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_366_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(366),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(107),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_365_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(365),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(106),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_364_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(364),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(105),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_363_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(363),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(104),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_362_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(362),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(103),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_361_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(361),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(102),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_360_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(360),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(101),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_359_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(359),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(100),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_358_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(358),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(99),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_357_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(357),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(98),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_356_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(356),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(97),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_355_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(355),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(96),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_354_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(354),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(95),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_353_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(353),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(94),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_352_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(352),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(93),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_351_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(351),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(92),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_350_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(350),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(91),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_349_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(349),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(90),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_348_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(348),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(89),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_347_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(347),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(88),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_346_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(346),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(87),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_345_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(345),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(86),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_344_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(344),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(85),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_343_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(343),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(84),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_342_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(342),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(83),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_341_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(341),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(82),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_340_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(340),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(81),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_339_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(339),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(80),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_338_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(338),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(79),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_337_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(337),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(78),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_336_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(336),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(77),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_335_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(335),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(76),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_334_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(334),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(75),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_333_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(333),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(74),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_332_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(332),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(73),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_331_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(331),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(72),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_330_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(330),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(71),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_329_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(329),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(70),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_328_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(328),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(69),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_327_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(327),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(68),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_326_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(326),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(67),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_325_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(325),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(66),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_324_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(324),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(65),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_323_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(323),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(64),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_322_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(322),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(63),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_321_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(321),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(62),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_320_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(320),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(61),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_319_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(319),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_319__G1\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_318_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(318),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_318__G1\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_317_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(317),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_317__G1\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_316_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(316),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_316__G1\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_315_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(315),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_314_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(314),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(55),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_313_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(313),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(54),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_312_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(312),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(53),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_311_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(311),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(52),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_310_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(310),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(51),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_309_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(309),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(50),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_308_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(308),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(49),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_307_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(307),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(48),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_306_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(306),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(47),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_305_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(305),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(46),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_304_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(304),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(45),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_303_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(303),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(44),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_302_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(302),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(43),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_301_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(301),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(42),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_300_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(300),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(41),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_299_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(299),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(40),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_298_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(298),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(39),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_297_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(297),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(38),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_296_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(296),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(37),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_295_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(295),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(36),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_294_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(294),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(35),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_293_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(293),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(34),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_292_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(292),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(33),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_291_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(291),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(32),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_290_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(290),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(31),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_289_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(289),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(30),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_288_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(288),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(29),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_287_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(287),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(28),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_286_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(286),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(27),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_285_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(285),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(26),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_284_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(284),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(25),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_283_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(283),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(24),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_282_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(282),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(23),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_281_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(281),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(22),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_280_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(280),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(21),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_279_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(279),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(20),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_278_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(278),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(19),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_277_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(277),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(18),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_276_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(276),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(17),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_275_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(275),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(16),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_274_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(274),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(15),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_273_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(273),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(14),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_272_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(272),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(13),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_271_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(271),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(12),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_270_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(270),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(11),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_269_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(269),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(10),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_268_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(268),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(9),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_267_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(267),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(8),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_266_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(266),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(7),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_265_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(265),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(6),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_264_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(264),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(5),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_263_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(263),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(4),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_262_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(262),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(3),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_261_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(261),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(2),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_260_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(260),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(1),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_259_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(259),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_8\(0),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_258_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(258),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_258__N_5_I\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4357\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_230_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(230),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF\(1),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_228_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(228),
d => \GRLFPC2_0.FPO.FRAC\(3),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_226_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(226),
d => \GRLFPC2_0.FPO.FRAC\(5),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_225_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(225),
d => \GRLFPC2_0.FPO.FRAC\(6),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_224_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(224),
d => \GRLFPC2_0.FPO.FRAC\(7),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_223_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(223),
d => \GRLFPC2_0.FPO.FRAC\(8),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_222_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(222),
d => \GRLFPC2_0.FPO.FRAC\(9),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_221_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(221),
d => \GRLFPC2_0.FPO.FRAC\(10),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_220_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(220),
d => \GRLFPC2_0.FPO.FRAC\(11),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_219_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(219),
d => \GRLFPC2_0.FPO.FRAC\(12),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_218_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(218),
d => \GRLFPC2_0.FPO.FRAC\(13),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_217_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(217),
d => \GRLFPC2_0.FPO.FRAC\(14),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_216_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(216),
d => \GRLFPC2_0.FPO.FRAC\(15),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_215_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(215),
d => \GRLFPC2_0.FPO.FRAC\(16),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_214_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(214),
d => \GRLFPC2_0.FPO.FRAC\(17),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_213_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(213),
d => \GRLFPC2_0.FPO.FRAC\(18),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_212_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(212),
d => \GRLFPC2_0.FPO.FRAC\(19),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_211_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(211),
d => \GRLFPC2_0.FPO.FRAC\(20),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_210_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(210),
d => \GRLFPC2_0.FPO.FRAC\(21),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_209_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(209),
d => \GRLFPC2_0.FPO.FRAC\(22),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_208_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(208),
d => \GRLFPC2_0.FPO.FRAC\(23),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_207_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(207),
d => \GRLFPC2_0.FPO.FRAC\(24),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_206_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(206),
d => \GRLFPC2_0.FPO.FRAC\(25),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_205_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(205),
d => \GRLFPC2_0.FPO.FRAC\(26),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_204_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(204),
d => \GRLFPC2_0.FPO.FRAC\(27),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_203_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(203),
d => \GRLFPC2_0.FPO.FRAC\(28),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_202_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(202),
d => N_27260,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27259,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
N_27258_I <= not N_27258;
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_201_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(201),
d => N_27262,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27261,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_200_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(200),
d => N_27264,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27263,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_199_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(199),
d => N_27266,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27265,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_198_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(198),
d => N_27268,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27267,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_197_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(197),
d => N_27270,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27269,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_196_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(196),
d => N_27272,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27271,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_195_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(195),
d => N_27274,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27273,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_194_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(194),
d => N_27276,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27275,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_193_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(193),
d => N_27278,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27277,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_192_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(192),
d => N_27280,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27279,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_191_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(191),
d => N_27282,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27281,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_190_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(190),
d => N_27284,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27283,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_189_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(189),
d => N_27286,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27285,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_188_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(188),
d => N_27288,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27287,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_187_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(187),
d => N_27290,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27289,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_186_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(186),
d => N_27292,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27291,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_185_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(185),
d => N_27294,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27293,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_184_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(184),
d => N_27296,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27295,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_183_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(183),
d => N_27298,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27297,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_182_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(182),
d => N_27300,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27299,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_181_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(181),
d => N_27302,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27301,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_180_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(180),
d => N_27304,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27303,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_179_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(179),
d => N_27306,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27305,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_178_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(178),
d => N_27308,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27307,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_177_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(177),
d => N_27310,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27309,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_176_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(176),
d => N_27312,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27311,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_175_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(175),
d => N_27314,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27313,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_174_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(174),
d => N_27316,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_231__G2\,
asdata => N_27315,
sload => N_27258_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_173_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(173),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(173),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_58_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(58),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_56_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10018\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10078\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_55_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10019\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10079\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_54_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10020\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10080\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_53_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10021\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10081\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_52_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10022\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10082\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_51_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10023\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_50_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10024\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10084\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_49_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10025\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10085\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_48_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10026\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10086\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_47_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10027\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10087\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_46_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10028\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10088\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_45_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10029\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10089\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_44_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10030\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10090\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_43_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10031\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10091\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_42_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10032\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10092\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_41_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10033\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10093\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_40_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10034\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10094\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_39_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10035\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10095\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_38_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10036\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10096\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_37_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10037\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10097\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_36_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10038\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10098\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_35_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10039\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10099\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_34_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10040\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10100\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_33_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10041\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10101\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_32_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10042\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10102\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_31_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10043\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10103\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_30_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10044\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10104\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_29_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10045\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10105\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_28_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10046\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10106\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_27_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10047\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10107\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_26_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10048\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10108\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_25_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10049\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10109\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_24_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10050\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10110\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_23_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10051\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10111\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_22_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10052\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10112\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_21_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10053\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10113\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_20_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10054\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10114\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_19_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10055\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10115\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_18_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10056\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10116\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
GRLFPC2_0_R_MK_HOLDN2: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.HOLDN2\,
d => \GRLFPC2_0.R.MK.HOLDN1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_RST2: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.RST2\,
d => \GRLFPC2_0.R.MK.RST_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_LDOP_RET: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.HOLDN_O\,
d => N_13,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_LDOP_RET_3: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.COMB.LOCKGEN.LOCKI_O_3\,
d => \GRLFPC2_0.N_3477_1_I\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_LDOP_RET_6: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O_3\(0),
d => N_14,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_RST_RET: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.COMB.ANNULFPU_1_O\,
d => \GRLFPC2_0.COMB.ANNULFPU_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_RST_RET_2: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.RST2_O\,
d => \GRLFPC2_0.R.MK.RST2\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_RST_RET_6: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.HOLDN2_O\,
d => \GRLFPC2_0.R.MK.HOLDN2\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_A_SEQERR_RET_3: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.N_1837_O\,
d => \GRLFPC2_0.N_76_I\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_I_PC_RET_60: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.V.I.EXEC_0_SQMUXA_O\,
d => N_37343_I_0,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_A_ST_RET: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.COMB.FPDECODE.ST_O\,
d => \GRLFPC2_0.COMB.FPDECODE.ST\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_A_AFQ_RET_5: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(0),
d => N_14,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_A_AFQ_RET_2: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.COMB.LOCKGEN.LOCKI_O\,
d => \GRLFPC2_0.N_3477_1_I\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_E_AFSR_RET: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.AFSR_O\,
d => \GRLFPC2_0.R.A.AFSR\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_E_AFQ_RET_1: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.N_1830_O\,
d => \GRLFPC2_0.N_1685\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_E_AFQ_RET: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.AFQ_O\,
d => \GRLFPC2_0.R.A.AFQ\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_M_AFSR_RET: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.E.AFSR_O\,
d => \GRLFPC2_0.R.M.AFSR_RET_0_0_G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_M_AFQ_RET_1: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.N_1829_O\,
d => \GRLFPC2_0.N_1683\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_M_AFQ_RET: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.E.AFQ_O\,
d => \GRLFPC2_0.R.M.AFQ_RET_0_0_G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_M_SEQERR: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.N_554\,
d => \GRLFPC2_0.N_553\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_E_SEQERR: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.N_553\,
d => \GRLFPC2_0.R.E.SEQERR_0_0_G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_A_RS2D: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RS2D\,
d => \GRLFPC2_0.COMB.RS2D_1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_A_RS1D: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RS1D\,
d => \GRLFPC2_0.COMB.RS1D_1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_X_RDD: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.X.RDD\,
d => \GRLFPC2_0.N_559\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_M_RDD: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.N_559\,
d => \GRLFPC2_0.N_558\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_E_RDD: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.N_558\,
d => \GRLFPC2_0.N_557\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_A_RDD: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.N_557\,
d => \GRLFPC2_0.R.A.RDD_0_0_G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_X_SEQERR: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.X.SEQERR\,
d => \GRLFPC2_0.N_554\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_A_LD: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.LD\,
d => \GRLFPC2_0.R.A.LD_0_0_G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_A_FPOP: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.FPOP\,
d => \GRLFPC2_0.R.A.FPOP_0_0_G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_I_EXEC: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.EXEC\,
d => N_37428,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_FTT_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.FTT\(2),
d => \GRLFPC2_0.R.FSR.FTT_0_0_2__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_FTT_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.FTT\(0),
d => \GRLFPC2_0.R.FSR.FTT_0_0_0__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_FSR_NONSTD: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.NONSTD\,
d => \GRLFPC2_0.R.FSR.NONSTD_0_0_G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_I_RDD: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RDD\,
d => N_37429,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_X_LD: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.X.LD\,
d => \GRLFPC2_0.R.X.LD_0_0_G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_X_FPOP: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.X.FPOP\,
d => \GRLFPC2_0.R.X.FPOP_0_0_G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_X_AFSR: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.X.AFSR\,
d => \GRLFPC2_0.R.X.AFSR_0_0_G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_X_AFQ: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.X.AFQ\,
d => \GRLFPC2_0.R.X.AFQ_0_0_G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_M_LD: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.M.LD\,
d => \GRLFPC2_0.R.M.LD_0_0_G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_M_FPOP: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.M.FPOP\,
d => \GRLFPC2_0.R.M.FPOP_0_0_G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_E_LD: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.E.LD\,
d => \GRLFPC2_0.R.E.LD_0_0_G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_E_FPOP: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.E.FPOP\,
d => \GRLFPC2_0.COMB.V.E.FPOP_1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_HOLDN1: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.HOLDN1\,
d => \GRLFPC2_0.N_2103\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_BUSY2_RET_1: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.BUSY_O\,
d => \GRLFPC2_0.N_2105\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
RST_I <= not N_11;
GRLFPC2_0_R_MK_BUSY2_RET: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.COMB.ANNULFPU_1_O_0\,
d => \GRLFPC2_0.COMB.ANNULFPU_1\,
clk => N_12,
clrn => VCC,
sclr => RST_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sload => GND);
GRLFPC2_0_R_MK_BUSY_RET_5: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.RST2_O_0\,
d => \GRLFPC2_0.R.MK.RST2\,
clk => N_12,
clrn => VCC,
sclr => RST_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sload => GND);
GRLFPC2_0_R_MK_BUSY_RET_4: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.RST_O_0\,
d => \GRLFPC2_0.N_2111\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_BUSY_RET_3: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.HOLDN2_O_0\,
d => \GRLFPC2_0.R.MK.HOLDN2\,
clk => N_12,
clrn => VCC,
sclr => RST_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sload => GND);
GRLFPC2_0_R_MK_BUSY_RET_2: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.HOLDN1_O_0\,
d => \GRLFPC2_0.R.MK.HOLDN1\,
clk => N_12,
clrn => VCC,
sclr => RST_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(0),
d => N_329,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(1),
d => N_330,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(2),
d => N_331,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(3),
d => N_332,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(4),
d => N_333,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_5_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(5),
d => N_334,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_6_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(6),
d => N_335,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_7_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(7),
d => N_336,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_8_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(8),
d => N_337,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_9_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(9),
d => N_338,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(10),
d => N_339,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_11_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(11),
d => N_340,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_12_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(12),
d => N_341,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_13_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(13),
d => N_342,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_14_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(14),
d => N_343,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(15),
d => N_344,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_16_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(16),
d => N_345,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_17_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(17),
d => N_346,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_18_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(18),
d => N_347,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_19_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(19),
d => N_348,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_20_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(20),
d => N_349,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_21_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(21),
d => N_350,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_22_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(22),
d => N_351,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_23_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(23),
d => N_352,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_24_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(24),
d => N_353,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_25_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(25),
d => N_354,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_26_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(26),
d => N_355,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_27_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(27),
d => N_356,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_28_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(28),
d => N_357,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_29_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(29),
d => N_358,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_30_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(30),
d => N_359,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_31_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(31),
d => N_360,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(0),
d => \GRLFPC2_0.R.E.STDATA_1_0_0__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(1),
d => \GRLFPC2_0.R.E.STDATA_1_0_1__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(2),
d => \GRLFPC2_0.R.E.STDATA_1_0_2__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(3),
d => \GRLFPC2_0.R.E.STDATA_1_0_3__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(4),
d => \GRLFPC2_0.R.E.STDATA_1_0_4__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_5_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(5),
d => \GRLFPC2_0.R.E.STDATA_1_0_5__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_6_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(6),
d => \GRLFPC2_0.R.E.STDATA_1_0_6__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_7_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(7),
d => \GRLFPC2_0.R.E.STDATA_1_0_7__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_8_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(8),
d => \GRLFPC2_0.R.E.STDATA_1_0_8__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_9_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(9),
d => \GRLFPC2_0.R.E.STDATA_1_0_9__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(10),
d => \GRLFPC2_0.R.E.STDATA_1_0_10__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_11_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(11),
d => \GRLFPC2_0.R.E.STDATA_1_0_11__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_12_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(12),
d => \GRLFPC2_0.R.E.STDATA_1_0_12__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_13_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(13),
d => \GRLFPC2_0.R.E.STDATA_1_0_13__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_14_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(14),
d => \GRLFPC2_0.R.E.STDATA_1_0_14__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(15),
d => \GRLFPC2_0.R.E.STDATA_1_0_15__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_16_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(16),
d => \GRLFPC2_0.R.E.STDATA_1_0_16__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_17_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(17),
d => \GRLFPC2_0.R.E.STDATA_1_0_17__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_18_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(18),
d => \GRLFPC2_0.R.E.STDATA_1_0_18__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_19_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(19),
d => \GRLFPC2_0.R.E.STDATA_1_0_19__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_20_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(20),
d => \GRLFPC2_0.R.E.STDATA_1_0_20__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_21_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(21),
d => \GRLFPC2_0.R.E.STDATA_1_0_21__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_22_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(22),
d => \GRLFPC2_0.R.E.STDATA_1_0_22__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_23_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(23),
d => \GRLFPC2_0.R.E.STDATA_1_0_23__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_24_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(24),
d => \GRLFPC2_0.R.E.STDATA_1_0_24__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_25_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(25),
d => \GRLFPC2_0.R.E.STDATA_1_0_25__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_26_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(26),
d => \GRLFPC2_0.R.E.STDATA_1_0_26__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_27_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(27),
d => \GRLFPC2_0.R.E.STDATA_1_0_27__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_28_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(28),
d => \GRLFPC2_0.R.E.STDATA_1_0_28__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_29_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(29),
d => \GRLFPC2_0.R.E.STDATA_1_0_29__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_30_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(30),
d => \GRLFPC2_0.R.E.STDATA_1_0_30__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_31_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(31),
d => \GRLFPC2_0.R.E.STDATA_1_0_31__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_RD_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.RD\(0),
d => \GRLFPC2_0.R.FSR.RD_0_0_0__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_RD_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.RD\(1),
d => \GRLFPC2_0.R.FSR.RD_0_0_1__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_TEM_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.TEM\(0),
d => \GRLFPC2_0.R.FSR.TEM_1_0_0__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_TEM_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.TEM\(1),
d => \GRLFPC2_0.R.FSR.TEM_1_0_1__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_TEM_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.TEM\(2),
d => \GRLFPC2_0.R.FSR.TEM_1_0_2__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_TEM_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.TEM\(3),
d => \GRLFPC2_0.R.FSR.TEM_1_0_3__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_TEM_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.TEM\(4),
d => \GRLFPC2_0.R.FSR.TEM_1_0_4__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_STATE_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.STATE\(0),
d => \GRLFPC2_0.R.STATE_0_0_0__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_STATE_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.STATE\(1),
d => \GRLFPC2_0.R.STATE_0_0_1__I0_I_1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RF1REN_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RF1REN\(2),
d => \GRLFPC2_0.N_3150\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RF1REN_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RF1REN\(1),
d => N_37431,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RF2REN_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RF2REN\(2),
d => N_37432,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RF2REN_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RF2REN\(1),
d => N_37433,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_FCC_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_CCZ(0),
d => \GRLFPC2_0.R.FSR.FCC_0_0_0__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_FCC_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_CCZ(1),
d => \GRLFPC2_0.R.FSR.FCC_0_0_1__G1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_AEXC_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.AEXC\(0),
d => \GRLFPC2_0.R.FSR.AEXC_1_0_0__I0_I_0\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_AEXC_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.AEXC\(1),
d => \GRLFPC2_0.R.FSR.AEXC_1_0_1__I0_I_1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_AEXC_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.AEXC\(2),
d => \GRLFPC2_0.R.FSR.AEXC_1_0_2__I0_I_0\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_AEXC_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.AEXC\(3),
d => \GRLFPC2_0.R.FSR.AEXC_1_0_3__I0_I_1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_AEXC_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.AEXC\(4),
d => \GRLFPC2_0.R.FSR.AEXC_1_0_4__I0_I_0\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_CEXC_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.CEXC\(0),
d => \GRLFPC2_0.R.FSR.CEXC_1_0_0__I0_I_1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_CEXC_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.CEXC\(1),
d => \GRLFPC2_0.R.FSR.CEXC_1_0_1__I0_I_0\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_CEXC_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.CEXC\(2),
d => \GRLFPC2_0.R.FSR.CEXC_1_0_2__I0_I_1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_CEXC_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.CEXC\(3),
d => \GRLFPC2_0.R.FSR.CEXC_1_0_3__I0_I_0\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_CEXC_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.CEXC\(4),
d => \GRLFPC2_0.R.FSR.CEXC_1_0_4__I0_I_1\,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_CC_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.CC\(0),
d => \GRLFPC2_0.R.I.CC_0_0_0__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_CC_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.CC\(1),
d => \GRLFPC2_0.R.I.CC_0_0_1__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_AFQ_RET_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(73),
d => N_87,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_AFQ_RET_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(74),
d => N_88,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_AFQ_RET_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(58),
d => N_72,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_AFQ_RET_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(59),
d => N_73,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_AFQ_RET_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(60),
d => N_74,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_AFQ_RET_5_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(61),
d => N_75,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_AFQ_RET_6_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(62),
d => N_76,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_AFQ_RET_7_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(63),
d => N_77,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_AFQ_RET_8_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(69),
d => N_83,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_AFQ_RET_9_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(70),
d => N_84,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_SEQERR_RET_4_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.STATE_O\(0),
d => \GRLFPC2_0.R.STATE\(0),
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_SEQERR_RET_4_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.STATE_O\(1),
d => \GRLFPC2_0.R.STATE\(1),
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(285),
d => N_299,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(286),
d => N_300,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(287),
d => N_301,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(288),
d => N_302,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(289),
d => N_303,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_5_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(290),
d => N_304,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_6_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(291),
d => N_305,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_7_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(292),
d => N_306,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_8_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(293),
d => N_307,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_9_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(294),
d => N_308,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(295),
d => N_309,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_11_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(296),
d => N_310,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_12_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(297),
d => N_311,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_13_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(298),
d => N_312,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_14_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(299),
d => N_313,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(300),
d => N_314,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_16_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(301),
d => N_315,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_17_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(302),
d => N_316,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_18_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(303),
d => N_317,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_19_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(304),
d => N_318,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_20_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(305),
d => N_319,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_21_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(306),
d => N_320,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_22_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(307),
d => N_321,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_23_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(308),
d => N_322,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_24_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(309),
d => N_323,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_25_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(310),
d => N_324,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_26_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(311),
d => N_325,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_27_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(312),
d => N_326,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_28_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(313),
d => N_327,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_29_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(314),
d => N_328,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(2),
d => \GRLFPC2_0.FPCI_O\(285),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(3),
d => \GRLFPC2_0.FPCI_O\(286),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(4),
d => \GRLFPC2_0.FPCI_O\(287),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(5),
d => \GRLFPC2_0.FPCI_O\(288),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(6),
d => \GRLFPC2_0.FPCI_O\(289),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_5_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(7),
d => \GRLFPC2_0.FPCI_O\(290),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_6_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(8),
d => \GRLFPC2_0.FPCI_O\(291),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_7_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(9),
d => \GRLFPC2_0.FPCI_O\(292),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_8_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(10),
d => \GRLFPC2_0.FPCI_O\(293),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_9_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(11),
d => \GRLFPC2_0.FPCI_O\(294),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(12),
d => \GRLFPC2_0.FPCI_O\(295),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_11_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(13),
d => \GRLFPC2_0.FPCI_O\(296),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_12_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(14),
d => \GRLFPC2_0.FPCI_O\(297),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_13_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(15),
d => \GRLFPC2_0.FPCI_O\(298),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_14_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(16),
d => \GRLFPC2_0.FPCI_O\(299),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(17),
d => \GRLFPC2_0.FPCI_O\(300),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_16_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(18),
d => \GRLFPC2_0.FPCI_O\(301),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_17_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(19),
d => \GRLFPC2_0.FPCI_O\(302),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_18_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(20),
d => \GRLFPC2_0.FPCI_O\(303),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_19_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(21),
d => \GRLFPC2_0.FPCI_O\(304),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_20_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(22),
d => \GRLFPC2_0.FPCI_O\(305),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_21_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(23),
d => \GRLFPC2_0.FPCI_O\(306),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_22_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(24),
d => \GRLFPC2_0.FPCI_O\(307),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_23_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(25),
d => \GRLFPC2_0.FPCI_O\(308),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_24_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(26),
d => \GRLFPC2_0.FPCI_O\(309),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_25_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(27),
d => \GRLFPC2_0.FPCI_O\(310),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_26_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(28),
d => \GRLFPC2_0.FPCI_O\(311),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_27_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(29),
d => \GRLFPC2_0.FPCI_O\(312),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_28_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(30),
d => \GRLFPC2_0.FPCI_O\(313),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_29_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_O\(31),
d => \GRLFPC2_0.FPCI_O\(314),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_9__G2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_MOV_RET_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(44),
d => N_58,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_MOV_RET_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(45),
d => N_59,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_MOV_RET_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(46),
d => N_60,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_MOV_RET_5_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(47),
d => N_61,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_MOV_RET_6_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(48),
d => N_62,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_MOV_RET_7_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(49),
d => N_63,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_MOV_RET_8_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(50),
d => N_64,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_MOV_RET_9_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(51),
d => N_65,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_MOV_RET_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O\(52),
d => N_66,
clk => N_12,
clrn => VCC,
ena => N_13,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_EXC_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.EXC\(0),
d => \GRLFPC2_0.R.I.EXC_MB\(0),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_EXC_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.EXC\(1),
d => \GRLFPC2_0.R.I.EXC_2_0_1__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_EXC_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.EXC\(2),
d => \GRLFPC2_0.R.I.EXC_2_0_2__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_EXC_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.EXC\(3),
d => \GRLFPC2_0.R.I.EXC_2_0_3__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_EXC_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.EXC\(4),
d => \GRLFPC2_0.R.I.EXC_2_0_4__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_1876_2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_MK_LDOP_RET_4_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.STATE_O_3\(0),
d => \GRLFPC2_0.R.STATE\(0),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_MK_LDOP_RET_4_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.STATE_O_3\(1),
d => \GRLFPC2_0.R.STATE\(1),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_MK_LDOP_RET_1_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O_3\(73),
d => N_87,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_MK_LDOP_RET_1_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O_3\(74),
d => N_88,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_MK_LDOP_RET_1_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O_0\(63),
d => N_77,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_MK_LDOP_RET_1_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O_0\(62),
d => N_76,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_MK_LDOP_RET_1_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O_0\(61),
d => N_75,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_MK_LDOP_RET_1_5_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O_0\(60),
d => N_74,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_MK_LDOP_RET_1_6_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O_0\(59),
d => N_73,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_MK_LDOP_RET_1_7_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O_0\(69),
d => N_83,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_MK_LDOP_RET_1_8_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPCI_O_0\(70),
d => N_84,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RS1_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RS1\(0),
d => \GRLFPC2_0.COMB.RS1_1\(0),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RS1_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RS1\(1),
d => \GRLFPC2_0.COMB.RS1_1\(1),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RS1_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RS1\(2),
d => \GRLFPC2_0.COMB.RS1_1\(2),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RS1_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RS1\(3),
d => \GRLFPC2_0.COMB.RS1_1\(3),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RS1_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RS1\(4),
d => \GRLFPC2_0.COMB.RS1_1\(4),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(0),
d => \GRLFPC2_0.FPO.FRAC\(3),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(1),
d => \GRLFPC2_0.FPO.FRAC\(4),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(2),
d => \GRLFPC2_0.FPO.FRAC\(5),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(3),
d => \GRLFPC2_0.FPO.FRAC\(6),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(4),
d => \GRLFPC2_0.FPO.FRAC\(7),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_5_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(5),
d => \GRLFPC2_0.FPO.FRAC\(8),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_6_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(6),
d => \GRLFPC2_0.FPO.FRAC\(9),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_7_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(7),
d => \GRLFPC2_0.FPO.FRAC\(10),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_8_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(8),
d => \GRLFPC2_0.FPO.FRAC\(11),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_9_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(9),
d => \GRLFPC2_0.FPO.FRAC\(12),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(10),
d => \GRLFPC2_0.FPO.FRAC\(13),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_11_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(11),
d => \GRLFPC2_0.FPO.FRAC\(14),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_12_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(12),
d => \GRLFPC2_0.FPO.FRAC\(15),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_13_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(13),
d => \GRLFPC2_0.FPO.FRAC\(16),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_14_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(14),
d => \GRLFPC2_0.FPO.FRAC\(17),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(15),
d => \GRLFPC2_0.FPO.FRAC\(18),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_16_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(16),
d => \GRLFPC2_0.FPO.FRAC\(19),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_17_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(17),
d => \GRLFPC2_0.FPO.FRAC\(20),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_18_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(18),
d => \GRLFPC2_0.FPO.FRAC\(21),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_19_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(19),
d => \GRLFPC2_0.FPO.FRAC\(22),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_20_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(20),
d => \GRLFPC2_0.FPO.FRAC\(23),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_21_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(21),
d => \GRLFPC2_0.FPO.FRAC\(24),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_22_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(22),
d => \GRLFPC2_0.FPO.FRAC\(25),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_23_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(23),
d => \GRLFPC2_0.FPO.FRAC\(26),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_24_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(24),
d => \GRLFPC2_0.FPO.FRAC\(27),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_25_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(25),
d => \GRLFPC2_0.FPO.FRAC\(28),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_26_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(26),
d => \GRLFPC2_0.FPO.FRAC\(29),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_27_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(27),
d => \GRLFPC2_0.FPO.FRAC\(30),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_28_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(28),
d => \GRLFPC2_0.FPO.FRAC\(31),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_60_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(60),
d => \GRLFPC2_0.FPO.EXP\(8),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_61_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(61),
d => \GRLFPC2_0.FPO.EXP\(9),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_62_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(62),
d => \GRLFPC2_0.FPO.EXP\(10),
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.N_54\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RS2_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RS2\(0),
d => \GRLFPC2_0.COMB.RS2_1\(0),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RS2_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RS2\(1),
d => \GRLFPC2_0.COMB.RS2_1\(1),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RS2_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RS2\(2),
d => \GRLFPC2_0.COMB.RS2_1\(2),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RS2_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RS2\(3),
d => \GRLFPC2_0.COMB.RS2_1\(3),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RS2_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RS2\(4),
d => \GRLFPC2_0.COMB.RS2_1\(4),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_RNI3OL9_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffff0fffff")
port map (
combout => N_61587_I_0,
dataf => \GRLFPC2_0.FPI.LDOP_1_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(5),
datad => \GRLFPC2_0.R.MK.RST2_0\,
datac => N_11);
GRLFPC2_0_FPI_LDOP_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff3000000")
port map (
combout => \GRLFPC2_0.FPI.LDOP_1_0\,
dataf => \GRLFPC2_0.R.MK.RST\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7920_I_A7_10\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7920_I_A7_6\,
datac => \GRLFPC2_0.R.STATE_O_3\(1),
datab => \GRLFPC2_0.R.STATE_O_3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_5_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(5),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_RST2_0: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.RST2_0\,
d => \GRLFPC2_0.R.MK.RST\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_FPI_LDOP_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff00ff")
port map (
combout => \GRLFPC2_0.FPI.LDOP_0\,
dataf => \GRLFPC2_0.FPI.LDOP_1_1\,
datae => \GRLFPC2_0.R.MK.RST2_1\,
datad => N_11);
GRLFPC2_0_FPI_LDOP_4: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff3000000")
port map (
combout => \GRLFPC2_0.FPI.LDOP_1_1\,
dataf => \GRLFPC2_0.R.MK.RST\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7920_I_A7_10\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7920_I_A7_6\,
datac => \GRLFPC2_0.R.STATE_O_3\(1),
datab => \GRLFPC2_0.R.STATE_O_3\(0));
GRLFPC2_0_R_MK_RST2_1: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.RST2_1\,
d => \GRLFPC2_0.R.MK.RST\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_RST_RET_0_RNIQF2I: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000f000000000")
port map (
combout => \GRLFPC2_0.R.MK.RST_0\,
dataf => \GRLFPC2_0.R.MK.RST_4_0\,
datae => \GRLFPC2_0.R.MK.RST2_2\,
datad => \GRLFPC2_0.R.MK.RST2_O_1\,
datac => \GRLFPC2_0.COMB.ANNULFPU_1_O_1\);
GRLFPC2_0_COMB_V_MK_RST_1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f000000000000000")
port map (
combout => \GRLFPC2_0.R.MK.RST_4_0\,
dataf => \GRLFPC2_0.R.MK.HOLDN2\,
datae => \GRLFPC2_0.HOLDN_O\,
datad => \GRLFPC2_0.FPO.BUSY_O\,
datac => \GRLFPC2_0.R.MK.HOLDN2_O\);
GRLFPC2_0_R_MK_RST2_2: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.RST2_2\,
d => \GRLFPC2_0.R.MK.RST\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_RST_RET_0: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.RST2_O_1\,
d => \GRLFPC2_0.R.MK.RST2\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_RST_RET_1: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.COMB.ANNULFPU_1_O_1\,
d => \GRLFPC2_0.COMB.ANNULFPU_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(0),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_1\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_RNO_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffa080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_3\,
datad => N_33794,
datac => N_29262_1,
datab => N_33795,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(0),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_RNO_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffa080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_3\,
datad => N_33794,
datac => N_29262_1,
datab => N_33795,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(0),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_5\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2_RNO_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffa080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_3\,
datad => N_33794,
datac => N_29262_1,
datab => N_33795,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(0),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_6\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3_RNO_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffa080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_3\,
datad => N_33794,
datac => N_29262_1,
datab => N_33795,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(0),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_7\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4_RNO_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffa080")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_3\,
datad => N_33794,
datac => N_29262_1,
datab => N_33795,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_17_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_1\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_RNO_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_10\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_12\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8714\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9349\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9373\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_17_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(17),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_3\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_RNO_17_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_10\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_12\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8714\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9349\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_9373\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_16_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI_0\(10),
clk => N_12,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_0_16_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI_0\(10),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_16__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_1: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_RETI_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNI6ERR_13_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"faf0fefcaa00eecc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_RETI_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(375),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(13));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_6: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_RETI_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_6_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"faf0fefcaa00eecc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_RETI_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(375),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIKDSA6_20_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f0f00000f0f0fd02")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datae => \GRLFPC2_0.FPI.LDOP_0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(20),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_1_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_1_RNO_10_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"f0f00000f0f0fd02")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datae => \GRLFPC2_0.FPI.LDOP_0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(20),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_RNO_0_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000fcf0fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(83),
dataf => N_65771_RETO,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_RNO_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO\,
dataa => CPI_D_INST_RETO(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"faffcafffa00ca00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10936_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN13_RESVEC_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(241));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000101ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10936_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10931\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7352\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM6\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_COMPUTECONST_UN13_RESVEC_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN13_RESVEC_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_31_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(31),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_32_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(32),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_29_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(29),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(29),
clk => N_12,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_241_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(241),
d => N_37418,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"faffcafffa00ca00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10936_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN13_RESVEC_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(241));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000101ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10936_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10931\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7352\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM6\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_COMPUTECONST_UN13_RESVEC_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN13_RESVEC_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_31_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(31),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_32_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(32),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_29_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(29),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(29),
clk => N_12,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1_241_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(241),
d => N_37418,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_RNI1FHI_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0f000fff0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_0\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_42_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(42),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_0\(15),
d => N_66970,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_43_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(43),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_RNI4FHI_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffff0f000fff0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(3),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_1\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_42_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(42),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_1_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_1\(15),
d => N_66970,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_43_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(43),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2_RNINTPE_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_2\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2_42_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(42),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_2_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_2\(15),
d => N_66970,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3_RNIPTPE_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_3\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3_42_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(42),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_3_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_3\(15),
d => N_66970,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4_RNIQTPE_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_4\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4_42_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(42),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_4_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_4\(15),
d => N_66970,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5_RNISTPE_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_1\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(1),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_5\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5_42_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(42),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_5_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_5\(15),
d => N_66970,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_2_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_2\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_56_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(56),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10018\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10078\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_24_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(24),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10050\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10110\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_3_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_3\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_54_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(54),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10020\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10080\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_22_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(22),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10052\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10112\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
GRLFPC2_0_FPI_LDOP_5: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff3000000")
port map (
combout => \GRLFPC2_0.FPI.LDOP_1_2\,
dataf => \GRLFPC2_0.R.MK.RST_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_I_A7_10_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_I_A7_6_0\,
datac => \GRLFPC2_0.R.STATE_O_3_0\(1),
datab => \GRLFPC2_0.R.STATE_O_3_0\(0));
GRLFPC2_0_FPI_LDOP_5_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000f000000000")
port map (
combout => \GRLFPC2_0.R.MK.RST_1\,
dataf => \GRLFPC2_0.R.MK.RST_4\,
datae => \GRLFPC2_0.R.MK.RST2\,
datad => \GRLFPC2_0.R.MK.RST2_O\,
datac => \GRLFPC2_0.COMB.ANNULFPU_1_O\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_232__G2_0_7920_I_A7\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0030000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_I_A7_10_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7920_I_A7_7\,
datae => \GRLFPC2_0.HOLDN_O\,
datad => \GRLFPC2_0.FPCI_O_0\(61),
datac => \GRLFPC2_0.FPCI_O_0\(62),
datab => \GRLFPC2_0.FPCI_O_0\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_232__G2_0_I_A7_0\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000f0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_I_A7_6_0\,
dataf => \GRLFPC2_0.FPCI_O_3\(0),
datae => \GRLFPC2_0.FPCI_O_0\(63),
datad => \GRLFPC2_0.FPCI_O_3\(73),
datac => \GRLFPC2_0.COMB.LOCKGEN.LOCKI_O_3\);
\GRLFPC2_0_R_MK_LDOP_RET_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.STATE_O_3_0\(1),
d => \GRLFPC2_0.R.STATE\(1),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_MK_LDOP_RET_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.STATE_O_3_0\(0),
d => \GRLFPC2_0.R.STATE\(0),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"5f0050005f305030")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19_0\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(244),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_NORMDETECT_NOTSLFROMNORM_19_0_A2_0_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0c0c0f0f0c0f0c0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19_0\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM12\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_244_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(244),
d => N_37415,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2_31_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(31),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2_32_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(32),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2_43_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(43),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_9: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC_RETI\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIGJ2IDT2_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffff0000f000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SM0_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_2_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0_N_5_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_1_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0_M3_I_A3_0_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_RNIE3QJME3_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"4c4c4c4444444c44")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_2_0\,
dataf => N_27316,
datae => N_27258,
datad => N_27315,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_RNIG14OGE3_0_68_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000f0f0f000f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0_N_5_0\,
dataf => N_27316,
datae => N_27258,
datad => N_27315,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_RNIPSLS5_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f3f0f3f0f3")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_1_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_49_I\,
datac => \GRLFPC2_0.FPI.LDOP_0_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIPHE9_0_3_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0fff0fff03f30")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0_M3_I_A3_0_0\,
dataf => \GRLFPC2_0.FPI.LDOP_1_2\,
datae => \GRLFPC2_0.R.MK.RST2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datab => N_11);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_4_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_4\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_55_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(55),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10019\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10079\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_23_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(23),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10051\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10111\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_5_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_5\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1_55_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(55),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10019\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10079\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1_23_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(23),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10051\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10111\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_1_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_6_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_6\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_2_55_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(55),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10019\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10079\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_2_23_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(23),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10051\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10111\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_7_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_7\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_53_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(53),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10021\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10081\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_21_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(21),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10053\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10113\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_8\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_8_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_8\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1_53_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(53),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10021\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10081\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1_21_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(21),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10053\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10113\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_1_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_9\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_9_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_9\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_2_53_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(53),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10021\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10081\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_2_21_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(21),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10053\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10113\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_10\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_10_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_10\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_25_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(25),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10049\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10109\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_57_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(57),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10017\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10077\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_1_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(8),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_11\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_11_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_11\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1_25_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(25),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10049\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10109\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1_57_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(57),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10017\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10077\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_2_8_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff0000ff00ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(8),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_12\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_12_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_12\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_2_25_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(25),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10049\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10109\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_2_57_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(57),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10017\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10077\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SS0_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff3fffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_2_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0_N_5_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_1_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0_M3_I_A3_0_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"4c4c4c4444444c44")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_2_1\,
dataf => N_27316,
datae => N_27258,
datad => N_27315,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SS0_0_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000f0f0f000f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0_N_5_1\,
dataf => N_27316,
datae => N_27258,
datad => N_27315,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"e0eee0ee00000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4897_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_1\,
datae => N_27258,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\,
datac => N_27315,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
datag => N_27316);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SS0_0_RNO_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f0f3f0f3f0f3")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_1_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_49_I\,
datac => \GRLFPC2_0.FPI.LDOP_0_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SS0_0_RNO_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fff0fff0fff03f30")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0_M3_I_A3_0_1\,
dataf => \GRLFPC2_0.FPI.LDOP_1_2\,
datae => \GRLFPC2_0.R.MK.RST2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datab => N_11);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN24_ZERO_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000f33")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5833_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_0\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_3\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_3\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_2_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_0\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_1_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_0\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_13_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_3_23_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_3\(23),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10051\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10111\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_3_55_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_3\(55),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10019\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10079\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN18_ZERO_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33ffffffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5828_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_1\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_4\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_4\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_3_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_1\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_2_5_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_1\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_14_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_4_23_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_4\(23),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10051\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10111\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_4_55_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_4\(55),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10019\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10079\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000fffeeefe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(2),
dataf => N_65516_0,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7778_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM12_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7777_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(31));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M14S2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM12_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7352\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_RNO_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_1\,
dataf => N_65496,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_0\,
datac => N_65775);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_YY_0_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"0000323200033232")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7778_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7352\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM6\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_XX_0_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000bbbbbbb8")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7777_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7350\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_SUB_0_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc0fffffcc0fff")
port map (
combout => N_65516_0,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3_31_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(31),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000fffeeefe")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
dataf => N_65516_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7778_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM12_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7777_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(31));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M14S2_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffffffffc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM12_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7352\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1_RNO_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000f0000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_2\,
dataf => N_65496,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_0\,
datac => N_65775);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_YY_1_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"0000323200033232")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7778_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7352\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM6\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_XX_1_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000bbbbbbb8")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7777_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7350\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_SUB_1_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00cc0fffffcc0fff")
port map (
combout => N_65516_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(2),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4_31_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(31),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0f0f0303030f03")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3632_0\,
dataf => N_27316,
datae => N_27258,
datad => N_27315,
datac => N_65549_0,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA_SUB_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffff00ffff0000")
port map (
combout => N_65549_0,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_I\,
datae => N_65719,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_0_68_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000000000c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4506_0\,
dataf => \GRLFPC2_0.FPI.LDOP_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(12),
datad => \GRLFPC2_0.R.MK.RST2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(47),
datab => N_11);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6_RNI0C6R_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"8888888888888880")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5105_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN12_SRTOSTICKY_1_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_6\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_6\(15));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN12_SRTOSTICKY: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN12_SRTOSTICKY_1_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(8),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6_42_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_6\(42),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_6_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_6\(15),
d => N_66970,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_RNIHOJ8_58_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00ff000000ff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_0\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(58),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_58_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(58),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(58),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_8_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(8),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_8__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_19_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(19),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_20_RNIOROM: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000ff00ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10800_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5346_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_12: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_RETI_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_18: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349_RETI\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_20: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5346_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5346_RETI\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_21_RNIUROM: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10743_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5346_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_21: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_0_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5365_RETI_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_26: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5349_RETI\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_27: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5346_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5346_RETI\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_32_RNIEPRJ3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f0000000d")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(84),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO_0\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_0\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_65_RNIG1E21: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333030033330000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO_0\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_TZ_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datab => CPI_D_INST_RETO(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_28_RNIJ1E21: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c333003300330033")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO_0\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(84));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_400_RNIBQ6O_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datae => N_65488_RETO_0,
datad => D_N_7_RETO_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_32: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_0\(1),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M\(1),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_33: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_38: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_50_RNIEPRJ3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f0000000d")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(84),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO_1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_65_RNIG1E21_7: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333030033330000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO_1\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_TZ_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datab => CPI_D_INST_RETO(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_28_RNIJ1E21_6: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c333003300330033")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO_1\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(84));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_400_RNIBQ6O_10: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datae => N_65488_RETO_0,
datad => D_N_7_RETO_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_50: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_1\(1),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M\(1),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_51: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_56: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_60_RNIDPRJ3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f0000000d")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(84),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO_2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO_2\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_65_RNIG1E21_6: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333030033330000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO_2\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_TZ_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datab => CPI_D_INST_RETO(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_28_RNIJ1E21_5: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c333003300330033")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO_2\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(84));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_400_RNIBQ6O_8: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datae => N_65488_RETO_0,
datad => D_N_7_RETO_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_60: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_2\(1),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M\(1),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_61: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO_2\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_62: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO_2\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_71_RNILPRJ3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f0000000d")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(84),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO_3\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO_3\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_3\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_65_RNIG1E21_4: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333030033330000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO_3\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_TZ_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datab => CPI_D_INST_RETO(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_28_RNIJ1E21_4: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c333003300330033")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO_3\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(84));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_400_RNIBQ6O_4: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datae => N_65488_RETO_0,
datad => D_N_7_RETO_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_63: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_3\(1),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M\(1),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_66: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO_3\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_71: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO_3\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_72_RNIOPRJ3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f0000000d")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(84),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO_4\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO_4\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_4\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO_4\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_65_RNIG1E21_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333030033330000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO_4\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_TZ_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datab => CPI_D_INST_RETO(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_28_RNIJ1E21_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c333003300330033")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO_4\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(84));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_400_RNIBQ6O_7: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datae => N_65488_RETO_0,
datad => D_N_7_RETO_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_72: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_4\(1),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M\(1),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_73: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO_4\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_76: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO_4\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_80_RNIUPRJ3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f0000000d")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(84),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO_5\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO_5\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_5\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO_5\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO_5\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_65_RNIG1E21_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333030033330000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO_5\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_TZ_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datab => CPI_D_INST_RETO(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_28_RNIJ1E21_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c333003300330033")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO_5\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(84));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_400_RNIBQ6O_6: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datae => N_65488_RETO_0,
datad => D_N_7_RETO_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_77: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_5\(1),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M\(1),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_79: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO_5\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_80: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO_5\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_81_RNIOPRJ3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f0000000d")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(84),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO_6\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO_6\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_6\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO_6\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO_6\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_65_RNIG1E21_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333030033330000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO_6\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_TZ_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datab => CPI_D_INST_RETO(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_28_RNIJ1E21_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c333003300330033")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO_6\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(84));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_400_RNIBQ6O_5: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datae => N_65488_RETO_0,
datad => D_N_7_RETO_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_81: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_6\(1),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M\(1),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_83: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO_6\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_84: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO_6\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_87_RNI9QRJ3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f0000000d")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(84),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO_7\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO_7\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_7\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO_7\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_65_RNIG1E21_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3333030033330000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO_7\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_TZ_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(65),
datab => CPI_D_INST_RETO(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_28_RNIJ1E21_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"c333003300330033")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO_7\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(84));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_400_RNIBQ6O_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datae => N_65488_RETO_0,
datad => D_N_7_RETO_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_87: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_7\(1),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M\(1),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_88: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO_7\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_99: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO_7\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_0_RNIJIIK_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000012003300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_248\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_0_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000300f300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(56));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_100: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_101: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_102: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_103: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_104: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(81),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_1_RNIF3JK_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000012003300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_249\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_1_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000300f300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(56));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_105: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_106: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_107: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_108: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_109: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(81),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_2_RNIU6KK_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000012003300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_250\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_2\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_2_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000300f300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_2\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(56));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_110: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_2\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_111: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_2\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_112: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_2\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_113: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_2\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_114: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_2\(81),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_3_RNIQNKK_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000012003300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_251\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_3\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_3_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000300f300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_3\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(56));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_115: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_3\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_116: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_3\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_117: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_3\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_118: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_3\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_119: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_3\(81),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_4_RNI9RLK_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000012003300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_4\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_4\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_4_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000300f300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_4\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(56));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_120: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_4\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_121: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_4\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_122: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_4\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_123: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_4\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_124: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_4\(81),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_5_RNI5CMK_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000012003300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_5\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_5\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_5\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_5_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000300f300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_5\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(56));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_125: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_5\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_126: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_5\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_127: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_5\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_128: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_5\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_129: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_5\(81),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_6_RNIKFNK_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000012003300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_6\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_6\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_6\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_6\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_6\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_6_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000300f300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_6\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(56));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_130: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_6\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_131: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_6\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_132: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_6\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_133: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_6\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_134: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_6\(81),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_8_RNIJGOK_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000012003300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_7\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_7\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_7\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_7\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_8_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000300f300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_7\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(56));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_135: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_7\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_136: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_7\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_137: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_7\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_138: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_7\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_139: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_7\(81),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_9_RNI2KPK_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000012003300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(81),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_8\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_8\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_8\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_8\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_8\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_0_A2_9_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000300f300")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1094_RETO_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(56));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_140: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_RETO_8\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_141: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0_RETO_8\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_2_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_142: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO_8\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_143: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102_RETO_8\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1102\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_144: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_8\(81),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_145_RNICGL32: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf000022230000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(85),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_8\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_0\,
dataa => CPI_D_INST_RETO_0(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_55_RNIR4BR_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff0fff0ccf0ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_0\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_400_RNIBQ6O_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_8\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datae => N_65488_RETO_0,
datad => D_N_7_RETO_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_145: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_146: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_147: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_148: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_0(10),
d => N_63,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_149_RNI1SL32: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf000022230000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(85),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_9\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_1\,
dataa => CPI_D_INST_RETO_1(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_55_RNIR4BR: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff0fff0ccf0ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_1\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_400_RNIBQ6O_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_9\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datae => N_65488_RETO_0,
datad => D_N_7_RETO_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_149: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_150: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_151: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_152: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_1(10),
d => N_63,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_153_RNI80M32: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf000022230000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(85),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_10\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_2\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_2\,
dataa => CPI_D_INST_RETO_2(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_55_RNIR4BR_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff0fff0ccf0ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_2\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_400_RNIBQ6O_15: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_10\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datae => N_65488_RETO_0,
datad => D_N_7_RETO_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_153: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_2\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_154: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_2\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_155: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_2\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_156: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_2(10),
d => N_63,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_157_RNIF4M32: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf000022230000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_274\(85),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_11\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_3\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_3\,
dataa => CPI_D_INST_RETO_3(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_55_RNIR4BR_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff0fff0ccf0ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_3\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_400_RNIBQ6O_18: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_11\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datae => N_65488_RETO_0,
datad => D_N_7_RETO_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_157: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_3\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_158: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_3\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_159: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_3\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_160: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_3(10),
d => N_63,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_161_RNI5GM32: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf000022230000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_275\(85),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_12\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_4\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_4\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_4\,
dataa => CPI_D_INST_RETO_4(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_55_RNIS4BR_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff0fff0ccf0ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_4\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_9\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_400_RNIBQ6O_17: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_12\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datae => N_65488_RETO_0,
datad => D_N_7_RETO_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_161: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_4\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_162: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_4\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_163: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_4\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_164: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_4(10),
d => N_63,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_165_RNILGM32: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf000022230000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_276\(85),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_13\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_5\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_5\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_5\,
dataa => CPI_D_INST_RETO_5(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_55_RNIS4BR: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff0fff0ccf0ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_5\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_9\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_400_RNIBQ6O_16: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_13\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datae => N_65488_RETO_0,
datad => D_N_7_RETO_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_165: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_5\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_166: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_5\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_167: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_5\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_168: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_5(10),
d => N_63,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_169_RNILA872: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf000022230000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_277\(85),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_14\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_6\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_6\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_6\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_6\,
dataa => CPI_D_INST_RETO_6(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_55_RNI7JSU_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff0fff0ccf0ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_6\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_9\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_400_RNIBQ6O_11: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_14\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datae => N_65488_RETO_0,
datad => D_N_7_RETO_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_169: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_6\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_170: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_6\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_171: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_6\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_172: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_6(10),
d => N_63,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_173_RNISE872: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf000022230000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_278\(85),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_15\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_7\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_7\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_7\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_7\,
dataa => CPI_D_INST_RETO_7(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_55_RNI7JSU_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff0fff0ccf0ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_7\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_9\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_400_RNIBQ6O_14: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_15\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datae => N_65488_RETO_0,
datad => D_N_7_RETO_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_173: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_7\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_174: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_7\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_175: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_7\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_176: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_7(10),
d => N_63,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_177_RNI3J872: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf000022230000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_279\(85),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_16\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_8\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_8\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_8\,
dataa => CPI_D_INST_RETO_8(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_55_RNI7JSU: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0ff0fff0ccf0ccf0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_8\(5),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_9\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_400_RNIBQ6O_13: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_16\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datae => N_65488_RETO_0,
datad => D_N_7_RETO_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_177: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_8\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_178: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_8\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_179: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_8\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_180: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_8(10),
d => N_63,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_181_RNISEAB2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_252\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_17\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_0\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_9\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_9\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_0\,
dataa => CPI_D_INST_RETO_0(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_74_RNIB3U21_4: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c3cff3caa3caa3c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_0\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO5_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_400_RNIBQ6O_12: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_17\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datae => N_65488_RETO_0,
datad => D_N_7_RETO_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_181: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_9\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_182: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_9\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_183: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_184: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_0(8),
d => N_61,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_185_RNICFAB2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_18\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_10\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_10\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_1\,
dataa => CPI_D_INST_RETO_1(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_74_RNIB3U21_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c3cff3caa3caa3c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_1\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO5_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_400_RNIBQ6O_9: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_18\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
datae => N_65488_RETO_0,
datad => D_N_7_RETO_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_185: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_10\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_186: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_10\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_187: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_188: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_1(8),
d => N_61,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_189_RNIVGBB2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_19\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_11\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_11\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_2\,
dataa => CPI_D_INST_RETO_2(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_74_RNIB3U21_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c3cff3caa3caa3c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_2\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO5_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_400_RNI9G7O_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_19\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO_0,
datad => D_N_7_RETO_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_189: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_11\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_190: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_11\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_191: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_2\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_192: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_2(8),
d => N_61,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_193_RNI6LBB2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_20\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_3\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_12\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_12\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_3\,
dataa => CPI_D_INST_RETO_3(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_74_RNIB3U21_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c3cff3caa3caa3c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_3\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO5_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_400_RNI9G7O_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_20\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO_0,
datad => D_N_7_RETO_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_193: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_12\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_194: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_12\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_195: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_3\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_196: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_3(8),
d => N_61,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_200_RNI4HAB2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_21\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_4\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_13\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_13\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_4\,
dataa => CPI_D_INST_RETO_4(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_74_RNIB3U21_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c3cff3caa3caa3c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_4\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO5_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_400_RNI9G7O: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_21\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO_0,
datad => D_N_7_RETO_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_197: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_13\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_198: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_13\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_199: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_4\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_200: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_4(8),
d => N_61,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_201_RNIV37B2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_22\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_5\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_14\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_14\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_5\,
dataa => CPI_D_INST_RETO_5(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_74_RNIC3U21: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c3cff3caa3caa3c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_5\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_9\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO5_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_400_RNI9G7O_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_22\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO_0,
datad => D_N_7_RETO_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_201: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_14\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_202: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_14\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_203: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_5\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_204: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_5(8),
d => N_61,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_205_RNIQIOE2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_23\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_6\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_15\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_15\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_6\,
dataa => CPI_D_INST_RETO_6(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_74_RNINHF61_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c3cff3caa3caa3c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_6\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_9\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO5_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_400_RNI9G7O_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_23\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO_0,
datad => D_N_7_RETO_0,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_205: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_15\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_206: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_15\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_207: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_6\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_208: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_6(8),
d => N_61,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_209_RNIVEI03: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_24\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_7\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_16\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_16\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_7\,
dataa => CPI_D_INST_RETO_7(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_74_RNINHF61_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c3cff3caa3caa3c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_7\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_9\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO5_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47_RNIP01A1_21: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_24\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO,
datad => D_N_7_RETO,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_209: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_16\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_210: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_16\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_211: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_7\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_212: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_7(8),
d => N_61,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_213_RNI6JI03: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_25\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_8\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_17\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_17\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_8\,
dataa => CPI_D_INST_RETO_8(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_74_RNINHF61: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c3cff3caa3caa3c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_8\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_9\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO5_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47_RNIP01A1_20: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_25\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO,
datad => D_N_7_RETO,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_213: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_17\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_214: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_17\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_215: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_8\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_216: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_8(8),
d => N_61,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_217_RNIDNI03: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(79),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_26\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_9\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_18\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_18\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_9\,
dataa => CPI_D_INST_RETO_9(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_74_RNINHF61_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"3c3cff3caa3caa3c")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_9\(3),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_9\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO5_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47_RNIP01A1_19: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_26\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO,
datad => D_N_7_RETO,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_217: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_18\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_218: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_18\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_219: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413_RETO_9\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_413\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_220: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_9(8),
d => N_61,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_221_RNIEJK43: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(78),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_27\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_0\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_19\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_19\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(84),
dataa => CPI_D_INST_RETO_0(12));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_24_RNI32HA1_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"3bffb1f5ce0ae4a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_0\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO5_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_8\,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47_RNIP01A1_18: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_27\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO,
datad => D_N_7_RETO,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_221: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_19\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_222: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_19\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_223: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(84),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_224: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_0(12),
d => N_65,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_225_RNIUJK43: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(78),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_28\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_1\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_20\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_20\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(84),
dataa => CPI_D_INST_RETO_1(12));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_24_RNI32HA1_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"3bffb1f5ce0ae4a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_1\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO5_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_8\,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47_RNIP01A1_17: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_28\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO,
datad => D_N_7_RETO,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_225: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_20\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_226: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_20\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_227: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(84),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_228: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_1(12),
d => N_65,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_229_RNIJVK43: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(78),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_29\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_2\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_21\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_21\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_2\(84),
dataa => CPI_D_INST_RETO_2(12));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_24_RNI32HA1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"3bffb1f5ce0ae4a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_2\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO5_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_8\,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47_RNIP01A1_16: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_29\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO,
datad => D_N_7_RETO,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_229: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_21\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_230: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_21\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_231: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_2\(84),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_232: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_2(12),
d => N_65,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_233_RNIQ3L43: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(78),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_30\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_3\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_22\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_22\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_3\(84),
dataa => CPI_D_INST_RETO_3(12));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_24_RNI32HA1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"3bffb1f5ce0ae4a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_3\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO5_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_8\,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47_RNIP01A1_15: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_30\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO,
datad => D_N_7_RETO,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_233: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_22\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_234: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_22\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_235: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_3\(84),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_236: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_3(12),
d => N_65,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_237_RNI28L43: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(78),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_31\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_4\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_23\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_23\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_4\(84),
dataa => CPI_D_INST_RETO_4(12));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_24_RNI42HA1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"3bffb1f5ce0ae4a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_4\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO5_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_9\,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47_RNIP01A1_14: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_31\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO,
datad => D_N_7_RETO,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_237: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_23\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_238: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_23\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_239: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_4\(84),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_240: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_4(12),
d => N_65,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_241_RNI22783: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(78),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_32\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_5\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_24\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_24\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_5\(84),
dataa => CPI_D_INST_RETO_5(12));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_24_RNIFG2E1_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"3bffb1f5ce0ae4a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_5\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO5_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_9\,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47_RNIP01A1_13: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_32\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO,
datad => D_N_7_RETO,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_241: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_24\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_242: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_24\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_243: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_5\(84),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_244: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_5(12),
d => N_65,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_245_RNII2783: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(78),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_33\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_6\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_25\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_25\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_6\(84),
dataa => CPI_D_INST_RETO_6(12));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_24_RNIFG2E1_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"3bffb1f5ce0ae4a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_6\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO5_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_9\,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47_RNIP01A1_12: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_33\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO,
datad => D_N_7_RETO,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_245: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_25\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_246: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_25\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_247: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_6\(84),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_248: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_6(12),
d => N_65,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_249_RNI7E783: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_264\(78),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_34\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_7\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_26\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_26\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_7\(84),
dataa => CPI_D_INST_RETO_7(12));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_24_RNIFG2E1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"3bffb1f5ce0ae4a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_7\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO5_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_9\,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47_RNIP01A1_11: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_34\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO,
datad => D_N_7_RETO,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_249: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_26\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_250: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_26\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_251: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_7\(84),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_252: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_7(12),
d => N_65,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_253_RNIEI783: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_265\(78),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_35\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_8\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_27\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_27\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_8\(84),
dataa => CPI_D_INST_RETO_8(12));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_24_RNIFG2E1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"3bffb1f5ce0ae4a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_8\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(78),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO5_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_9\,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47_RNIP01A1_10: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_35\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO,
datad => D_N_7_RETO,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_253: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_27\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_254: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_27\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_255: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_8\(84),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_256: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_8(12),
d => N_65,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_257_RNI68M43: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_253\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_36\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_28\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_28\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(79),
dataa => CPI_D_INST_RETO_0(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_30_RNI02HA1_4: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"3bffb1f5ce0ae4a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_0\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_8\,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47_RNIP01A1_9: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_36\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO,
datad => D_N_7_RETO,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_257: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_28\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_258: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_28\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_259: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_0\(79),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_260: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_0(5),
d => N_58,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_261_RNIRJM43: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_254\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_37\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_29\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_29\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(79),
dataa => CPI_D_INST_RETO_1(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_30_RNI02HA1_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"3bffb1f5ce0ae4a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_1\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_8\,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47_RNIP01A1_8: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_37\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO,
datad => D_N_7_RETO,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_261: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_29\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_262: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_29\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_263: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_1\(79),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_264: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_1(5),
d => N_58,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_265_RNIBKM43: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_255\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_38\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_30\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_30\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_2\(79),
dataa => CPI_D_INST_RETO_2(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_30_RNI02HA1_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"3bffb1f5ce0ae4a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_2\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_8\,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47_RNIP01A1_7: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_38\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO,
datad => D_N_7_RETO,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_265: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_30\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_266: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_30\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_267: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_2\(79),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_268: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_2(5),
d => N_58,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_269_RNI00N43: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_256\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_39\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_3\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_31\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_31\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_3\(79),
dataa => CPI_D_INST_RETO_3(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_30_RNI02HA1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"3bffb1f5ce0ae4a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_3\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_8\,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47_RNIP01A1_6: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_39\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO,
datad => D_N_7_RETO,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_269: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_31\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_270: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_31\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_271: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_3\(79),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_272: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_3(5),
d => N_58,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_273_RNI74N43: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_257\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_40\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_4\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_32\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_32\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_4\(79),
dataa => CPI_D_INST_RETO_4(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_30_RNI02HA1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"3bffb1f5ce0ae4a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_4\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_8\,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47_RNIP01A1_5: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_40\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO,
datad => D_N_7_RETO,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_273: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_32\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_274: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_32\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_275: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_4\(79),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_276: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_4(5),
d => N_58,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_277_RNIF8N43: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_258\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_41\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_5\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_33\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_33\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_5\(79),
dataa => CPI_D_INST_RETO_5(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_30_RNI12HA1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"3bffb1f5ce0ae4a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_5\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_9\,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47_RNIP01A1_4: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_41\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO,
datad => D_N_7_RETO,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_277: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_33\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_278: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_33\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_279: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_5\(79),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_280: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_5(5),
d => N_58,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_281_RNIF2983: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_259\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_42\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_6\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_34\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_34\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_6\(79),
dataa => CPI_D_INST_RETO_6(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_30_RNICG2E1_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"3bffb1f5ce0ae4a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_6\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_9\,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47_RNIP01A1_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_42\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO,
datad => D_N_7_RETO,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_281: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_34\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_282: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_34\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_283: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_6\(79),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_284: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_6(5),
d => N_58,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_285_RNIV2983: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_43\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_7\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_35\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_35\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_7\(79),
dataa => CPI_D_INST_RETO_7(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_30_RNICG2E1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"3bffb1f5ce0ae4a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_7\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_9\,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47_RNIP01A1_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_43\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO,
datad => D_N_7_RETO,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_285: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_35\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_286: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_35\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_287: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_7\(79),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_288: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_7(5),
d => N_58,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_289_RNIKE983: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_261\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_44\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_8\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_36\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_36\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_8\(79),
dataa => CPI_D_INST_RETO_8(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_30_RNICG2E1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"3bffb1f5ce0ae4a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_8\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_9\,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47_RNIP01A1_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_44\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO,
datad => D_N_7_RETO,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_289: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_36\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_290: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_36\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_291: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_8\(79),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_292: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_8(5),
d => N_58,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_293_RNIRI983: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_262\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_45\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_9\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_37\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_37\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_9\(79),
dataa => CPI_D_INST_RETO_9(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_30_RNICG2E1_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"3bffb1f5ce0ae4a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_9\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_9\,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47_RNIP01A1_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_45\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO,
datad => D_N_7_RETO,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_293: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_37\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_294: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_37\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_295: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_9\(79),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_296: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_9(5),
d => N_58,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_300_RNIPE883: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf0000888c0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_263\(80),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_46\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_10\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_38\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_38\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_10\(79),
dataa => CPI_D_INST_RETO_10(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_30_RNICG2E1_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "on",
    lut_mask => X"3bffb1f5ce0ae4a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_10\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(80),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_1_CO3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_9\,
datag => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47_RNIP01A1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffefffefffefbfaf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_46\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO\,
datae => N_65488_RETO,
datad => D_N_7_RETO,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_297: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_38\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_298: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_38\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_299: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO_10\(79),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_300: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_10(5),
d => N_58,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_301_RNIEBDE1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000fcf0fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_266\(83),
dataf => N_65771_RETO_0,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_90_RNI0RBU_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fff00ff00ff00ff")
port map (
combout => N_65771_RETO_0,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO\,
datad => N_65609_RETO,
datac => CPI_D_INST_RETO(7));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_301: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_302: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_303: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_304: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_305_RNIUBDE1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000fcf0fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_267\(83),
dataf => N_65771_RETO_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_90_RNI0RBU_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fff00ff00ff00ff")
port map (
combout => N_65771_RETO_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO\,
datad => N_65609_RETO,
datac => CPI_D_INST_RETO(7));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_305: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_306: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_307: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_308: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_309_RNIJNDE1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000fcf0fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_268\(83),
dataf => N_65771_RETO_2,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_90_RNI0RBU_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fff00ff00ff00ff")
port map (
combout => N_65771_RETO_2,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO\,
datad => N_65609_RETO,
datac => CPI_D_INST_RETO(7));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_309: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO_2\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_310: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_2\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_311: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO_2\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_312: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO_2\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_313_RNIQRDE1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000fcf0fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_269\(83),
dataf => N_65771_RETO_3,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_90_RNI0RBU_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fff00ff00ff00ff")
port map (
combout => N_65771_RETO_3,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO\,
datad => N_65609_RETO,
datac => CPI_D_INST_RETO(7));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_313: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO_3\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_314: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_3\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_315: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO_3\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_316: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO_3\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_317_RNI10EE1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000fcf0fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_270\(83),
dataf => N_65771_RETO_4,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO_4\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO_4\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_90_RNI0RBU_7: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fff00ff00ff00ff")
port map (
combout => N_65771_RETO_4,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO\,
datad => N_65609_RETO,
datac => CPI_D_INST_RETO(7));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_317: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO_4\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_318: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_4\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_319: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO_4\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_320: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO_4\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_321_RNIMBEE1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000fcf0fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_271\(83),
dataf => N_65771_RETO_5,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO_5\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO_5\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_90_RNI0RBU_6: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fff00ff00ff00ff")
port map (
combout => N_65771_RETO_5,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO\,
datad => N_65609_RETO,
datac => CPI_D_INST_RETO(7));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_321: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO_5\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_322: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_5\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_323: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO_5\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_324: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO_5\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_325_RNI6CEE1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000fcf0fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272\(83),
dataf => N_65771_RETO_6,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO_6\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_6\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO_6\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO_6\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_90_RNI0RBU_5: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fff00ff00ff00ff")
port map (
combout => N_65771_RETO_6,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO\,
datad => N_65609_RETO,
datac => CPI_D_INST_RETO(7));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_325: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO_6\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_326: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_6\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_327: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO_6\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_328: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO_6\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_329_RNIRNEE1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000fcf0fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_273\(83),
dataf => N_65771_RETO_7,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO_7\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_7\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO_7\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO_7\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_90_RNI0RBU_4: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0fff00ff00ff00ff")
port map (
combout => N_65771_RETO_7,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO\,
datad => N_65609_RETO,
datac => CPI_D_INST_RETO(7));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_329: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_RETO_7\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_330: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_7\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_331: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6_RETO_7\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_6\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_332: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4_RETO_7\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_REST_N_4\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_333_RNIPH4O: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffff8fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_235\(82),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_0\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_0\,
dataa => CPI_D_INST_RETO_0(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_333: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_334: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_335: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_0\(3),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M\(3),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_336: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_337: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_338: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_0(11),
d => N_64,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_339_RNIG55O: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffff8fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_236\(82),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_1\,
dataa => CPI_D_INST_RETO_1(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_339: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_340: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_341: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_1\(3),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M\(3),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_342: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_343: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_344: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_1(11),
d => N_64,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_345_RNI2E5O: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffff8fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_237\(82),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_2\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_2\,
dataa => CPI_D_INST_RETO_2(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_345: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_2\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_346: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_2\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_347: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_2\(3),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M\(3),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_348: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_2\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_349: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_2\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_350: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_2(11),
d => N_64,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_351_RNIP16O: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffff8fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_238\(82),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_3\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_3\,
dataa => CPI_D_INST_RETO_3(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_351: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_3\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_352: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_3\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_353: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_3\(3),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M\(3),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_354: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_3\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_355: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_3\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_356: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_3(11),
d => N_64,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_357_RNI2E6O: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffff8fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_239\(82),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_4\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_4\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_4\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_4\,
dataa => CPI_D_INST_RETO_4(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_357: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_4\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_358: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_4\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_359: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_4\(3),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M\(3),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_360: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_4\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_361: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_4\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_362: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_4(11),
d => N_64,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_363_RNIBQ6O: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffff8fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_240\(82),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_5\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_5\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_5\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_5\,
dataa => CPI_D_INST_RETO_5(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_363: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_5\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_364: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_5\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_365: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_5\(3),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M\(3),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_366: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_5\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_367: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_5\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_368: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_5(11),
d => N_64,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_369_RNI2E7O: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffff8fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_241\(82),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_6\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_6\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_6\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_6\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_6\,
dataa => CPI_D_INST_RETO_6(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_369: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_6\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_370: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_6\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_371: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_6\(3),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M\(3),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_372: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_6\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_373: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_6\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_374: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_6(11),
d => N_64,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_375_RNIKM7O: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffff8fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_242\(82),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_7\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_7\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_7\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_7\,
dataa => CPI_D_INST_RETO_7(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_375: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_7\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_376: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_7\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_377: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_7\(3),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M\(3),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_378: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_7\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_379: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_7\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_380: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_7(11),
d => N_64,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_381_RNIBA8O: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffff8fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_243\(82),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_8\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_8\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_8\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_8\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_8\,
dataa => CPI_D_INST_RETO_8(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_381: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_8\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_382: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_8\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_383: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_8\(3),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M\(3),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_384: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_8\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_385: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_8\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_386: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_8(11),
d => N_64,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_387_RNIKM8O: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffffff8fff0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_244\(82),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_9\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_9\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_9\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_9\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_9\,
dataa => CPI_D_INST_RETO_9(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_387: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2_RETO_9\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G2\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_388: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D_RETO_9\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_D\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_389: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M_RETO_9\(3),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_M\(3),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_390: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1_RETO_9\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_391: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C_RETO_9\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_C\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_392: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO_9(11),
d => N_64,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN5_ZERO_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"33ff5f5fffccfafa")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_6163_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_0\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_3\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_5\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_5\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_3\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_1_7_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_0\(7),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_2\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_15_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_2\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_3_25_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_3\(25),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10049\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10109\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_5_55_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_5\(55),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10019\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10079\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_5_23_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_5\(23),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10051\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10111\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_3_57_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_3\(57),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10017\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10077\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
GRLFPC2_0_FPI_LDOP_6: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff00ff")
port map (
combout => \GRLFPC2_0.FPI.LDOP_0_0\,
dataf => \GRLFPC2_0.FPI.LDOP_1_1_0\,
datae => \GRLFPC2_0.R.MK.RST2_1_0\,
datad => N_11);
GRLFPC2_0_FPI_LDOP_7: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff3000000")
port map (
combout => \GRLFPC2_0.FPI.LDOP_1_1_0\,
dataf => \GRLFPC2_0.R.MK.RST\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7920_I_A7_10\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7920_I_A7_6\,
datac => \GRLFPC2_0.R.STATE_O_3\(1),
datab => \GRLFPC2_0.R.STATE_O_3\(0));
GRLFPC2_0_R_MK_RST2_3: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.RST2_1_0\,
d => \GRLFPC2_0.R.MK.RST\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_FPI_LDOP_8: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffff00ff")
port map (
combout => \GRLFPC2_0.FPI.LDOP_0_1\,
dataf => \GRLFPC2_0.FPI.LDOP_1_1_1\,
datae => \GRLFPC2_0.R.MK.RST2_1_1\,
datad => N_11);
GRLFPC2_0_FPI_LDOP_9: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff3000000")
port map (
combout => \GRLFPC2_0.FPI.LDOP_1_1_1\,
dataf => \GRLFPC2_0.R.MK.RST\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7920_I_A7_10\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7920_I_A7_6\,
datac => \GRLFPC2_0.R.STATE_O_3\(1),
datab => \GRLFPC2_0.R.STATE_O_3\(0));
GRLFPC2_0_R_MK_RST2_4: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.RST2_1_1\,
d => \GRLFPC2_0.R.MK.RST\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_393: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_8\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_393_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffcccf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_394: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_RETO_9\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_1\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_394_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffffffcccf")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_673_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_395: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_RETO_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_PCTRL_NEW_1_S_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000300000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_S_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_513\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_877_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_551\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_396: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_RETO_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_2\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CHECKOVANDDENORM_UN13_NOTPOSSIBLEOV_2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"8000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_2\,
dataf => \GRLFPC2_0.FPO.FRAC\(54),
datae => \GRLFPC2_0.FPO.FRAC\(52),
datad => \GRLFPC2_0.FPO.FRAC\(53),
datac => \GRLFPC2_0.FPO.FRAC\(49),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_397: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => N_65488_RETO_0,
d => N_65488_0,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_397_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0035ffffffffffff")
port map (
combout => N_65488_0,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_D\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0_0\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0\(9),
datac => N_27258,
datab => N_27310,
dataa => N_27309);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_398: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => D_N_7_RETO_0,
d => D_N_7_0,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_398_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000200010003")
port map (
combout => D_N_7_0,
dataf => N_44787,
datae => N_53932,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_663\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK\,
dataa => N_44786);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_399: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_RETO_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_I_O2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffa000ffffeccc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_399_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1846\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1539\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_411\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1852\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1839\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1618\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_400: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_RETO_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_M2_E_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_401: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_RETO_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_I_48: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff00f0fffff0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_I_0_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_475\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(67),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(66));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000000000000ffff")
port map (
combout => N_32738_1_0,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260_0\(84),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272_0\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_RNO_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000f0000000d")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_260_0\(84),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_I_M_RETO_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_RETO_0\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_IV_M_RETO_0\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_70_RETO_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1854_RETO_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_RNO_0_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"aaaf000022230000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_272_0\(85),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_61_RETO_9\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_0_1_RETO_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_RETO_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_RETO_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO_1\,
dataa => CPI_D_INST_RETO_1(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7_RNIVTPE_42_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000ff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_0\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE\(0),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_7\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_7\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7_42_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_7\(42),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_7_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_7\(15),
d => N_66970,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_13\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_16_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_13\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_51_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(51),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10023\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_19_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(19),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10055\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10115\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_1\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_14\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_17_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_14\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1_51_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(51),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10023\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1_19_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(19),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10055\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10115\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_1_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_15\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_18_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_15\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_2_51_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(51),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10023\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10083\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_2_19_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_2\(19),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10055\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10115\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffafcfaff0a0c0a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_0\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10934_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(243));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0d0c0c0c0d0c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10934_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7786\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM12\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10931\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_402: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC_RETI\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3_32_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(32),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5_31_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_5\(31),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2_29_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2\(29),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(29),
clk => N_12,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_243_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(243),
d => N_37416,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffafcfaff0a0c0a0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10934_1\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_6\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(243));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_4_1_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0f0d0c0c0c0d0c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10934_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7786\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_SM12\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10931\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_403: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC_2\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC_RETI\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4_32_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_4\(32),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6_31_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_6\(31),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3_29_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_3\(29),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(29),
clk => N_12,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1_243_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(243),
d => N_37416,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_0_A2: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000300000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_879_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_513_0\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_479_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(65));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_0_A2_RNO: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffffffffcccc00c0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1544\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1852\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1503\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1633\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1618\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_2_I_O2_0_83_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f3f3f3f3f3333333")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_513_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_458\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_426\,
datad => N_32738_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(67),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(66));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_0_O2_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f0fffffff0fff0f")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_479_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(71),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(74),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_65_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(65),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW_2\(65),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTABORTNULLEXC_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ff00ffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(75),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN39_ZERO_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000f33")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7065_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_2\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(20),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_4_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_2\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_2_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_0\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_13\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_19_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_3\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_20_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(20),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10054\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10114\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_52_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(52),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10022\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10082\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN33_ZERO_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0f33ffffffffffff")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_7057_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_3\(4),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(20),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_5_4_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_3\(4),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_7\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_3_2_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff00ffff0000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_1\(2),
dataf => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_13\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_0\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_20_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.UN1_GRFPULITE0_0_4\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4460_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1_20_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(20),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10054\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10114\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1_52_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH_1\(52),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10022\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4118\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10082\,
sload => N_61587_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_0_0_TZ_0_RNIM1VI843: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000004010101050")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_0\,
dataf => D_N_7_1,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_3\,
datad => N_65488_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_TZ_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(65));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CHECKOVANDDENORM_UN13_NOTPOSSIBLEOV_3: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"8000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_3\,
dataf => \GRLFPC2_0.FPO.FRAC\(54),
datae => \GRLFPC2_0.FPO.FRAC\(52),
datad => \GRLFPC2_0.FPO.FRAC\(53),
datac => \GRLFPC2_0.FPO.FRAC\(49),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN18_LOCOV_RNI2D3459_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0035ffffffffffff")
port map (
combout => N_65488_1,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_D\(7),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0_0\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0\(9),
datac => N_27258,
datab => N_27310,
dataa => N_27309);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_27_D_D_0_RNIQUBP2R2_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000200010003")
port map (
combout => D_N_7_1,
dataf => N_44787,
datae => N_53932,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_663\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK\,
dataa => N_44786);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_0_0_TZ_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"cc00cc00fff0ff00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0_0_TZ_0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1855\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_513\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_877_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_551\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_M2_E_1: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000000c00")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_N_3_1\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1856\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_3895\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN6_FEEDBACK\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_65_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_1\(65),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW_2\(65),
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_RNI27AB_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000000000f00000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_10075_0\,
dataf => \GRLFPC2_0.FPI.LDOP_1_3\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(6),
datad => \GRLFPC2_0.R.MK.RST2_3\,
datac => N_11);
GRLFPC2_0_FPI_LDOP_10: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"fffffffff3000000")
port map (
combout => \GRLFPC2_0.FPI.LDOP_1_3\,
dataf => \GRLFPC2_0.R.MK.RST\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7920_I_A7_10\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_232__G2_0_7920_I_A7_6\,
datac => \GRLFPC2_0.R.STATE_O_3\(1),
datab => \GRLFPC2_0.R.STATE_O_3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_6_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(6),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2\,
clk => N_12,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__N_5\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_RST2_5: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.RST2_3\,
d => \GRLFPC2_0.R.MK.RST_0\,
clk => N_12,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_V_STATE_2_SQMUXA0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000f000f000f000")
port map (
combout => \GRLFPC2_0.V.STATE_2_SQMUXA0\,
dataf => \GRLFPC2_0.R.I.EXC\(2),
datae => \GRLFPC2_0.R.FSR.TEM\(2),
datad => \GRLFPC2_0.COMB.UN1_MEXC_0\,
datac => \GRLFPC2_0.COMB.UN1_MEXC_1\);
GRLFPC2_0_V_STATE_2_SQMUXA: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff13ff130000ff13")
port map (
combout => \GRLFPC2_0.N_1495\,
dataf => \GRLFPC2_0.V.STATE_2_SQMUXA0\,
datae => \GRLFPC2_0.COMB.V.STATE12_0\,
datad => \GRLFPC2_0.N_1105\,
datac => \GRLFPC2_0.R.X.AFQ\,
datab => \GRLFPC2_0.R.X.SEQERR\,
dataa => \GRLFPC2_0.N_76_I\);
GRLFPC2_0_COMB_UN1_V_STATE0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ff00ff0000ff0000")
port map (
combout => \GRLFPC2_0.COMB.UN1_V.STATE0\,
dataf => \GRLFPC2_0.R.X.SEQERR\,
datae => \GRLFPC2_0.R.X.AFQ\,
datad => \GRLFPC2_0.N_1105\);
GRLFPC2_0_COMB_V_FSR_FCC80: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0fff0ff00f0f0ff")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.FCC80\,
dataf => \GRLFPC2_0.R.STATE\(0),
datae => \GRLFPC2_0.R.X.SEQERR\,
datad => \GRLFPC2_0.N_76_I\,
datac => \GRLFPC2_0.COMB.UN1_V.STATE0\);
GRLFPC2_0_COMB_V_FSR_FCC8: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"0000c00000000000")
port map (
combout => \GRLFPC2_0.N_1133\,
dataf => \GRLFPC2_0.COMB.V.FSR.FCC80\,
datae => \GRLFPC2_0.R.STATE\(0),
datad => \GRLFPC2_0.V.STATE_2_SQMUXA0\,
datac => \GRLFPC2_0.COMB.V.STATE12_0\,
datab => \GRLFPC2_0.COMB.ISFPOP2_1\);
GRLFPC2_0_V_FSR_CEXC_2_SQMUXA0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"00000000ffff0000")
port map (
combout => \GRLFPC2_0.V.FSR.CEXC_2_SQMUXA0\,
dataf => \GRLFPC2_0.N_1517\,
datae => \GRLFPC2_0.N_1171\);
GRLFPC2_0_V_FSR_CEXC_2_SQMUXA: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"d4fff4ff44444444")
port map (
combout => \GRLFPC2_0.V.FSR.CEXC_2_SQMUXA\,
dataf => \GRLFPC2_0.V.FSR.CEXC_2_SQMUXA0\,
datae => \GRLFPC2_0.COMB.ISFPOP2_1\,
datad => \GRLFPC2_0.COMB.V.STATE12_0\,
datac => \GRLFPC2_0.V.STATE_2_SQMUXA0\,
datab => \GRLFPC2_0.R.STATE\(0),
dataa => \GRLFPC2_0.COMB.V.FSR.FCC80\);
GRLFPC2_0_COMB_UN1_V_STATE0_0: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"000f00ff0000000f")
port map (
combout => \GRLFPC2_0.COMB.UN1_V.STATE0_0\,
dataf => \GRLFPC2_0.COMB.UN1_V.STATE0\,
datae => \GRLFPC2_0.R.X.SEQERR\,
datad => \GRLFPC2_0.R.STATE\(0),
datac => \GRLFPC2_0.R.STATE\(1));
GRLFPC2_0_COMB_UN1_V_STATE: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"7f55555500000000")
port map (
combout => N_37318_1,
dataf => \GRLFPC2_0.COMB.UN1_V.STATE0_0\,
datae => \GRLFPC2_0.COMB.UN1_MEXC_1\,
datad => \GRLFPC2_0.COMB.UN1_MEXC_0\,
datac => \GRLFPC2_0.R.FSR.TEM\(2),
datab => \GRLFPC2_0.R.I.EXC\(2),
dataa => \GRLFPC2_0.COMB.V.STATE12_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_00_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"f0fff0f0000ff0f0")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_00\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_0_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ccccccc333cc33cc")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN21_EXPXBUS\(0),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_00\,
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(43),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS0_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"ffff000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS0\,
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(10),
datae => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_6_\: stratixiii_lcell_comb generic map (
    shared_arith => "off",
    extended_lut => "off",
    lut_mask => X"d5f5d55580a08000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(6),
dataf => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS0\,
datae => RFO2_DATA1_RETO(3),
datad => \GRLFPC2_0.FPI.LDOP_I_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_4462_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(109),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0\(17));
N_11 <= RST_INTERNAL;
N_12 <= CLK_INTERNAL;
N_13 <= HOLDN_INTERNAL;
N_14 <= CPI_FLUSH_INTERNAL;
N_15 <= CPI_EXACK_INTERNAL;
N_16 <= CPI_A_RS1_INTERNAL;
N_17 <= CPI_A_RS1_INTERNAL_0;
N_18 <= CPI_A_RS1_INTERNAL_1;
N_19 <= CPI_A_RS1_INTERNAL_2;
N_20 <= CPI_A_RS1_INTERNAL_3;
N_21 <= CPI_D_PC_INTERNAL;
N_22 <= CPI_D_PC_INTERNAL_0;
N_23 <= CPI_D_PC_INTERNAL_1;
N_24 <= CPI_D_PC_INTERNAL_2;
N_25 <= CPI_D_PC_INTERNAL_3;
N_26 <= CPI_D_PC_INTERNAL_4;
N_27 <= CPI_D_PC_INTERNAL_5;
N_28 <= CPI_D_PC_INTERNAL_6;
N_29 <= CPI_D_PC_INTERNAL_7;
N_30 <= CPI_D_PC_INTERNAL_8;
N_31 <= CPI_D_PC_INTERNAL_9;
N_32 <= CPI_D_PC_INTERNAL_10;
N_33 <= CPI_D_PC_INTERNAL_11;
N_34 <= CPI_D_PC_INTERNAL_12;
N_35 <= CPI_D_PC_INTERNAL_13;
N_36 <= CPI_D_PC_INTERNAL_14;
N_37 <= CPI_D_PC_INTERNAL_15;
N_38 <= CPI_D_PC_INTERNAL_16;
N_39 <= CPI_D_PC_INTERNAL_17;
N_40 <= CPI_D_PC_INTERNAL_18;
N_41 <= CPI_D_PC_INTERNAL_19;
N_42 <= CPI_D_PC_INTERNAL_20;
N_43 <= CPI_D_PC_INTERNAL_21;
N_44 <= CPI_D_PC_INTERNAL_22;
N_45 <= CPI_D_PC_INTERNAL_23;
N_46 <= CPI_D_PC_INTERNAL_24;
N_47 <= CPI_D_PC_INTERNAL_25;
N_48 <= CPI_D_PC_INTERNAL_26;
N_49 <= CPI_D_PC_INTERNAL_27;
N_50 <= CPI_D_PC_INTERNAL_28;
N_51 <= CPI_D_PC_INTERNAL_29;
N_52 <= CPI_D_PC_INTERNAL_30;
N_53 <= CPI_D_INST_INTERNAL;
N_54 <= CPI_D_INST_INTERNAL_0;
N_55 <= CPI_D_INST_INTERNAL_1;
N_56 <= CPI_D_INST_INTERNAL_2;
N_57 <= CPI_D_INST_INTERNAL_3;
N_58 <= CPI_D_INST_INTERNAL_4;
N_59 <= CPI_D_INST_INTERNAL_5;
N_60 <= CPI_D_INST_INTERNAL_6;
N_61 <= CPI_D_INST_INTERNAL_7;
N_62 <= CPI_D_INST_INTERNAL_8;
N_63 <= CPI_D_INST_INTERNAL_9;
N_64 <= CPI_D_INST_INTERNAL_10;
N_65 <= CPI_D_INST_INTERNAL_11;
N_66 <= CPI_D_INST_INTERNAL_12;
N_67 <= CPI_D_INST_INTERNAL_13;
N_68 <= CPI_D_INST_INTERNAL_14;
N_69 <= CPI_D_INST_INTERNAL_15;
N_70 <= CPI_D_INST_INTERNAL_16;
N_71 <= CPI_D_INST_INTERNAL_17;
N_72 <= CPI_D_INST_INTERNAL_18;
N_73 <= CPI_D_INST_INTERNAL_19;
N_74 <= CPI_D_INST_INTERNAL_20;
N_75 <= CPI_D_INST_INTERNAL_21;
N_76 <= CPI_D_INST_INTERNAL_22;
N_77 <= CPI_D_INST_INTERNAL_23;
N_78 <= CPI_D_INST_INTERNAL_24;
N_79 <= CPI_D_INST_INTERNAL_25;
N_80 <= CPI_D_INST_INTERNAL_26;
N_81 <= CPI_D_INST_INTERNAL_27;
N_82 <= CPI_D_INST_INTERNAL_28;
N_83 <= CPI_D_INST_INTERNAL_29;
N_84 <= CPI_D_INST_INTERNAL_30;
N_85 <= CPI_D_CNT_INTERNAL;
N_86 <= CPI_D_CNT_INTERNAL_0;
N_87 <= CPI_D_TRAP_INTERNAL;
N_88 <= CPI_D_ANNUL_INTERNAL;
N_89 <= CPI_D_PV_INTERNAL;
N_90 <= CPI_A_PC_INTERNAL;
N_91 <= CPI_A_PC_INTERNAL_0;
N_92 <= CPI_A_PC_INTERNAL_1;
N_93 <= CPI_A_PC_INTERNAL_2;
N_94 <= CPI_A_PC_INTERNAL_3;
N_95 <= CPI_A_PC_INTERNAL_4;
N_96 <= CPI_A_PC_INTERNAL_5;
N_97 <= CPI_A_PC_INTERNAL_6;
N_98 <= CPI_A_PC_INTERNAL_7;
N_99 <= CPI_A_PC_INTERNAL_8;
N_100 <= CPI_A_PC_INTERNAL_9;
N_101 <= CPI_A_PC_INTERNAL_10;
N_102 <= CPI_A_PC_INTERNAL_11;
N_103 <= CPI_A_PC_INTERNAL_12;
N_104 <= CPI_A_PC_INTERNAL_13;
N_105 <= CPI_A_PC_INTERNAL_14;
N_106 <= CPI_A_PC_INTERNAL_15;
N_107 <= CPI_A_PC_INTERNAL_16;
N_108 <= CPI_A_PC_INTERNAL_17;
N_109 <= CPI_A_PC_INTERNAL_18;
N_110 <= CPI_A_PC_INTERNAL_19;
N_111 <= CPI_A_PC_INTERNAL_20;
N_112 <= CPI_A_PC_INTERNAL_21;
N_113 <= CPI_A_PC_INTERNAL_22;
N_114 <= CPI_A_PC_INTERNAL_23;
N_115 <= CPI_A_PC_INTERNAL_24;
N_116 <= CPI_A_PC_INTERNAL_25;
N_117 <= CPI_A_PC_INTERNAL_26;
N_118 <= CPI_A_PC_INTERNAL_27;
N_119 <= CPI_A_PC_INTERNAL_28;
N_120 <= CPI_A_PC_INTERNAL_29;
N_121 <= CPI_A_PC_INTERNAL_30;
N_122 <= CPI_A_INST_INTERNAL;
N_123 <= CPI_A_INST_INTERNAL_0;
N_124 <= CPI_A_INST_INTERNAL_1;
N_125 <= CPI_A_INST_INTERNAL_2;
N_126 <= CPI_A_INST_INTERNAL_3;
N_127 <= CPI_A_INST_INTERNAL_4;
N_128 <= CPI_A_INST_INTERNAL_5;
N_129 <= CPI_A_INST_INTERNAL_6;
N_130 <= CPI_A_INST_INTERNAL_7;
N_131 <= CPI_A_INST_INTERNAL_8;
N_132 <= CPI_A_INST_INTERNAL_9;
N_133 <= CPI_A_INST_INTERNAL_10;
N_134 <= CPI_A_INST_INTERNAL_11;
N_135 <= CPI_A_INST_INTERNAL_12;
N_136 <= CPI_A_INST_INTERNAL_13;
N_137 <= CPI_A_INST_INTERNAL_14;
N_138 <= CPI_A_INST_INTERNAL_15;
N_139 <= CPI_A_INST_INTERNAL_16;
N_140 <= CPI_A_INST_INTERNAL_17;
N_141 <= CPI_A_INST_INTERNAL_18;
N_142 <= CPI_A_INST_INTERNAL_19;
N_143 <= CPI_A_INST_INTERNAL_20;
N_144 <= CPI_A_INST_INTERNAL_21;
N_145 <= CPI_A_INST_INTERNAL_22;
N_146 <= CPI_A_INST_INTERNAL_23;
N_147 <= CPI_A_INST_INTERNAL_24;
N_148 <= CPI_A_INST_INTERNAL_25;
N_149 <= CPI_A_INST_INTERNAL_26;
N_150 <= CPI_A_INST_INTERNAL_27;
N_151 <= CPI_A_INST_INTERNAL_28;
N_152 <= CPI_A_INST_INTERNAL_29;
N_153 <= CPI_A_INST_INTERNAL_30;
N_154 <= CPI_A_CNT_INTERNAL;
N_155 <= CPI_A_CNT_INTERNAL_0;
N_156 <= CPI_A_TRAP_INTERNAL;
N_157 <= CPI_A_ANNUL_INTERNAL;
N_158 <= CPI_A_PV_INTERNAL;
N_159 <= CPI_E_PC_INTERNAL;
N_160 <= CPI_E_PC_INTERNAL_0;
N_161 <= CPI_E_PC_INTERNAL_1;
N_162 <= CPI_E_PC_INTERNAL_2;
N_163 <= CPI_E_PC_INTERNAL_3;
N_164 <= CPI_E_PC_INTERNAL_4;
N_165 <= CPI_E_PC_INTERNAL_5;
N_166 <= CPI_E_PC_INTERNAL_6;
N_167 <= CPI_E_PC_INTERNAL_7;
N_168 <= CPI_E_PC_INTERNAL_8;
N_169 <= CPI_E_PC_INTERNAL_9;
N_170 <= CPI_E_PC_INTERNAL_10;
N_171 <= CPI_E_PC_INTERNAL_11;
N_172 <= CPI_E_PC_INTERNAL_12;
N_173 <= CPI_E_PC_INTERNAL_13;
N_174 <= CPI_E_PC_INTERNAL_14;
N_175 <= CPI_E_PC_INTERNAL_15;
N_176 <= CPI_E_PC_INTERNAL_16;
N_177 <= CPI_E_PC_INTERNAL_17;
N_178 <= CPI_E_PC_INTERNAL_18;
N_179 <= CPI_E_PC_INTERNAL_19;
N_180 <= CPI_E_PC_INTERNAL_20;
N_181 <= CPI_E_PC_INTERNAL_21;
N_182 <= CPI_E_PC_INTERNAL_22;
N_183 <= CPI_E_PC_INTERNAL_23;
N_184 <= CPI_E_PC_INTERNAL_24;
N_185 <= CPI_E_PC_INTERNAL_25;
N_186 <= CPI_E_PC_INTERNAL_26;
N_187 <= CPI_E_PC_INTERNAL_27;
N_188 <= CPI_E_PC_INTERNAL_28;
N_189 <= CPI_E_PC_INTERNAL_29;
N_190 <= CPI_E_PC_INTERNAL_30;
N_191 <= CPI_E_INST_INTERNAL;
N_192 <= CPI_E_INST_INTERNAL_0;
N_193 <= CPI_E_INST_INTERNAL_1;
N_194 <= CPI_E_INST_INTERNAL_2;
N_195 <= CPI_E_INST_INTERNAL_3;
N_196 <= CPI_E_INST_INTERNAL_4;
N_197 <= CPI_E_INST_INTERNAL_5;
N_198 <= CPI_E_INST_INTERNAL_6;
N_199 <= CPI_E_INST_INTERNAL_7;
N_200 <= CPI_E_INST_INTERNAL_8;
N_201 <= CPI_E_INST_INTERNAL_9;
N_202 <= CPI_E_INST_INTERNAL_10;
N_203 <= CPI_E_INST_INTERNAL_11;
N_204 <= CPI_E_INST_INTERNAL_12;
N_205 <= CPI_E_INST_INTERNAL_13;
N_206 <= CPI_E_INST_INTERNAL_14;
N_207 <= CPI_E_INST_INTERNAL_15;
N_208 <= CPI_E_INST_INTERNAL_16;
N_209 <= CPI_E_INST_INTERNAL_17;
N_210 <= CPI_E_INST_INTERNAL_18;
N_211 <= CPI_E_INST_INTERNAL_19;
N_212 <= CPI_E_INST_INTERNAL_20;
N_213 <= CPI_E_INST_INTERNAL_21;
N_214 <= CPI_E_INST_INTERNAL_22;
N_215 <= CPI_E_INST_INTERNAL_23;
N_216 <= CPI_E_INST_INTERNAL_24;
N_217 <= CPI_E_INST_INTERNAL_25;
N_218 <= CPI_E_INST_INTERNAL_26;
N_219 <= CPI_E_INST_INTERNAL_27;
N_220 <= CPI_E_INST_INTERNAL_28;
N_221 <= CPI_E_INST_INTERNAL_29;
N_222 <= CPI_E_INST_INTERNAL_30;
N_223 <= CPI_E_CNT_INTERNAL;
N_224 <= CPI_E_CNT_INTERNAL_0;
N_225 <= CPI_E_TRAP_INTERNAL;
N_226 <= CPI_E_ANNUL_INTERNAL;
N_227 <= CPI_E_PV_INTERNAL;
N_228 <= CPI_M_PC_INTERNAL;
N_229 <= CPI_M_PC_INTERNAL_0;
N_230 <= CPI_M_PC_INTERNAL_1;
N_231 <= CPI_M_PC_INTERNAL_2;
N_232 <= CPI_M_PC_INTERNAL_3;
N_233 <= CPI_M_PC_INTERNAL_4;
N_234 <= CPI_M_PC_INTERNAL_5;
N_235 <= CPI_M_PC_INTERNAL_6;
N_236 <= CPI_M_PC_INTERNAL_7;
N_237 <= CPI_M_PC_INTERNAL_8;
N_238 <= CPI_M_PC_INTERNAL_9;
N_239 <= CPI_M_PC_INTERNAL_10;
N_240 <= CPI_M_PC_INTERNAL_11;
N_241 <= CPI_M_PC_INTERNAL_12;
N_242 <= CPI_M_PC_INTERNAL_13;
N_243 <= CPI_M_PC_INTERNAL_14;
N_244 <= CPI_M_PC_INTERNAL_15;
N_245 <= CPI_M_PC_INTERNAL_16;
N_246 <= CPI_M_PC_INTERNAL_17;
N_247 <= CPI_M_PC_INTERNAL_18;
N_248 <= CPI_M_PC_INTERNAL_19;
N_249 <= CPI_M_PC_INTERNAL_20;
N_250 <= CPI_M_PC_INTERNAL_21;
N_251 <= CPI_M_PC_INTERNAL_22;
N_252 <= CPI_M_PC_INTERNAL_23;
N_253 <= CPI_M_PC_INTERNAL_24;
N_254 <= CPI_M_PC_INTERNAL_25;
N_255 <= CPI_M_PC_INTERNAL_26;
N_256 <= CPI_M_PC_INTERNAL_27;
N_257 <= CPI_M_PC_INTERNAL_28;
N_258 <= CPI_M_PC_INTERNAL_29;
N_259 <= CPI_M_PC_INTERNAL_30;
N_260 <= CPI_M_INST_INTERNAL;
N_261 <= CPI_M_INST_INTERNAL_0;
N_262 <= CPI_M_INST_INTERNAL_1;
N_263 <= CPI_M_INST_INTERNAL_2;
N_264 <= CPI_M_INST_INTERNAL_3;
N_265 <= CPI_M_INST_INTERNAL_4;
N_266 <= CPI_M_INST_INTERNAL_5;
N_267 <= CPI_M_INST_INTERNAL_6;
N_268 <= CPI_M_INST_INTERNAL_7;
N_269 <= CPI_M_INST_INTERNAL_8;
N_270 <= CPI_M_INST_INTERNAL_9;
N_271 <= CPI_M_INST_INTERNAL_10;
N_272 <= CPI_M_INST_INTERNAL_11;
N_273 <= CPI_M_INST_INTERNAL_12;
N_274 <= CPI_M_INST_INTERNAL_13;
N_275 <= CPI_M_INST_INTERNAL_14;
N_276 <= CPI_M_INST_INTERNAL_15;
N_277 <= CPI_M_INST_INTERNAL_16;
N_278 <= CPI_M_INST_INTERNAL_17;
N_279 <= CPI_M_INST_INTERNAL_18;
N_280 <= CPI_M_INST_INTERNAL_19;
N_281 <= CPI_M_INST_INTERNAL_20;
N_282 <= CPI_M_INST_INTERNAL_21;
N_283 <= CPI_M_INST_INTERNAL_22;
N_284 <= CPI_M_INST_INTERNAL_23;
N_285 <= CPI_M_INST_INTERNAL_24;
N_286 <= CPI_M_INST_INTERNAL_25;
N_287 <= CPI_M_INST_INTERNAL_26;
N_288 <= CPI_M_INST_INTERNAL_27;
N_289 <= CPI_M_INST_INTERNAL_28;
N_290 <= CPI_M_INST_INTERNAL_29;
N_291 <= CPI_M_INST_INTERNAL_30;
N_292 <= CPI_M_CNT_INTERNAL;
N_293 <= CPI_M_CNT_INTERNAL_0;
N_294 <= CPI_M_TRAP_INTERNAL;
N_295 <= CPI_M_ANNUL_INTERNAL;
N_296 <= CPI_M_PV_INTERNAL;
N_297 <= CPI_X_PC_INTERNAL;
N_298 <= CPI_X_PC_INTERNAL_0;
N_299 <= CPI_X_PC_INTERNAL_1;
N_300 <= CPI_X_PC_INTERNAL_2;
N_301 <= CPI_X_PC_INTERNAL_3;
N_302 <= CPI_X_PC_INTERNAL_4;
N_303 <= CPI_X_PC_INTERNAL_5;
N_304 <= CPI_X_PC_INTERNAL_6;
N_305 <= CPI_X_PC_INTERNAL_7;
N_306 <= CPI_X_PC_INTERNAL_8;
N_307 <= CPI_X_PC_INTERNAL_9;
N_308 <= CPI_X_PC_INTERNAL_10;
N_309 <= CPI_X_PC_INTERNAL_11;
N_310 <= CPI_X_PC_INTERNAL_12;
N_311 <= CPI_X_PC_INTERNAL_13;
N_312 <= CPI_X_PC_INTERNAL_14;
N_313 <= CPI_X_PC_INTERNAL_15;
N_314 <= CPI_X_PC_INTERNAL_16;
N_315 <= CPI_X_PC_INTERNAL_17;
N_316 <= CPI_X_PC_INTERNAL_18;
N_317 <= CPI_X_PC_INTERNAL_19;
N_318 <= CPI_X_PC_INTERNAL_20;
N_319 <= CPI_X_PC_INTERNAL_21;
N_320 <= CPI_X_PC_INTERNAL_22;
N_321 <= CPI_X_PC_INTERNAL_23;
N_322 <= CPI_X_PC_INTERNAL_24;
N_323 <= CPI_X_PC_INTERNAL_25;
N_324 <= CPI_X_PC_INTERNAL_26;
N_325 <= CPI_X_PC_INTERNAL_27;
N_326 <= CPI_X_PC_INTERNAL_28;
N_327 <= CPI_X_PC_INTERNAL_29;
N_328 <= CPI_X_PC_INTERNAL_30;
N_329 <= CPI_X_INST_INTERNAL;
N_330 <= CPI_X_INST_INTERNAL_0;
N_331 <= CPI_X_INST_INTERNAL_1;
N_332 <= CPI_X_INST_INTERNAL_2;
N_333 <= CPI_X_INST_INTERNAL_3;
N_334 <= CPI_X_INST_INTERNAL_4;
N_335 <= CPI_X_INST_INTERNAL_5;
N_336 <= CPI_X_INST_INTERNAL_6;
N_337 <= CPI_X_INST_INTERNAL_7;
N_338 <= CPI_X_INST_INTERNAL_8;
N_339 <= CPI_X_INST_INTERNAL_9;
N_340 <= CPI_X_INST_INTERNAL_10;
N_341 <= CPI_X_INST_INTERNAL_11;
N_342 <= CPI_X_INST_INTERNAL_12;
N_343 <= CPI_X_INST_INTERNAL_13;
N_344 <= CPI_X_INST_INTERNAL_14;
N_345 <= CPI_X_INST_INTERNAL_15;
N_346 <= CPI_X_INST_INTERNAL_16;
N_347 <= CPI_X_INST_INTERNAL_17;
N_348 <= CPI_X_INST_INTERNAL_18;
N_349 <= CPI_X_INST_INTERNAL_19;
N_350 <= CPI_X_INST_INTERNAL_20;
N_351 <= CPI_X_INST_INTERNAL_21;
N_352 <= CPI_X_INST_INTERNAL_22;
N_353 <= CPI_X_INST_INTERNAL_23;
N_354 <= CPI_X_INST_INTERNAL_24;
N_355 <= CPI_X_INST_INTERNAL_25;
N_356 <= CPI_X_INST_INTERNAL_26;
N_357 <= CPI_X_INST_INTERNAL_27;
N_358 <= CPI_X_INST_INTERNAL_28;
N_359 <= CPI_X_INST_INTERNAL_29;
N_360 <= CPI_X_INST_INTERNAL_30;
N_361 <= CPI_X_CNT_INTERNAL;
N_362 <= CPI_X_CNT_INTERNAL_0;
N_363 <= CPI_X_TRAP_INTERNAL;
N_364 <= CPI_X_ANNUL_INTERNAL;
N_365 <= CPI_X_PV_INTERNAL;
N_366 <= CPI_LDDATA_INTERNAL;
N_367 <= CPI_LDDATA_INTERNAL_0;
N_368 <= CPI_LDDATA_INTERNAL_1;
N_369 <= CPI_LDDATA_INTERNAL_2;
N_370 <= CPI_LDDATA_INTERNAL_3;
N_371 <= CPI_LDDATA_INTERNAL_4;
N_372 <= CPI_LDDATA_INTERNAL_5;
N_373 <= CPI_LDDATA_INTERNAL_6;
N_374 <= CPI_LDDATA_INTERNAL_7;
N_375 <= CPI_LDDATA_INTERNAL_8;
N_376 <= CPI_LDDATA_INTERNAL_9;
N_377 <= CPI_LDDATA_INTERNAL_10;
N_378 <= CPI_LDDATA_INTERNAL_11;
N_379 <= CPI_LDDATA_INTERNAL_12;
N_380 <= CPI_LDDATA_INTERNAL_13;
N_381 <= CPI_LDDATA_INTERNAL_14;
N_382 <= CPI_LDDATA_INTERNAL_15;
N_383 <= CPI_LDDATA_INTERNAL_16;
N_384 <= CPI_LDDATA_INTERNAL_17;
N_385 <= CPI_LDDATA_INTERNAL_18;
N_386 <= CPI_LDDATA_INTERNAL_19;
N_387 <= CPI_LDDATA_INTERNAL_20;
N_388 <= CPI_LDDATA_INTERNAL_21;
N_389 <= CPI_LDDATA_INTERNAL_22;
N_390 <= CPI_LDDATA_INTERNAL_23;
N_391 <= CPI_LDDATA_INTERNAL_24;
N_392 <= CPI_LDDATA_INTERNAL_25;
N_393 <= CPI_LDDATA_INTERNAL_26;
N_394 <= CPI_LDDATA_INTERNAL_27;
N_395 <= CPI_LDDATA_INTERNAL_28;
N_396 <= CPI_LDDATA_INTERNAL_29;
N_397 <= CPI_LDDATA_INTERNAL_30;
N_398 <= CPI_DBG_ENABLE_INTERNAL;
N_399 <= CPI_DBG_WRITE_INTERNAL;
N_400 <= CPI_DBG_FSR_INTERNAL;
N_401 <= CPI_DBG_ADDR_INTERNAL;
N_402 <= CPI_DBG_ADDR_INTERNAL_0;
N_403 <= CPI_DBG_ADDR_INTERNAL_1;
N_404 <= CPI_DBG_ADDR_INTERNAL_2;
N_405 <= CPI_DBG_ADDR_INTERNAL_3;
N_406 <= CPI_DBG_DATA_INTERNAL;
N_407 <= CPI_DBG_DATA_INTERNAL_0;
N_408 <= CPI_DBG_DATA_INTERNAL_1;
N_409 <= CPI_DBG_DATA_INTERNAL_2;
N_410 <= CPI_DBG_DATA_INTERNAL_3;
N_411 <= CPI_DBG_DATA_INTERNAL_4;
N_412 <= CPI_DBG_DATA_INTERNAL_5;
N_413 <= CPI_DBG_DATA_INTERNAL_6;
N_414 <= CPI_DBG_DATA_INTERNAL_7;
N_415 <= CPI_DBG_DATA_INTERNAL_8;
N_416 <= CPI_DBG_DATA_INTERNAL_9;
N_417 <= CPI_DBG_DATA_INTERNAL_10;
N_418 <= CPI_DBG_DATA_INTERNAL_11;
N_419 <= CPI_DBG_DATA_INTERNAL_12;
N_420 <= CPI_DBG_DATA_INTERNAL_13;
N_421 <= CPI_DBG_DATA_INTERNAL_14;
N_422 <= CPI_DBG_DATA_INTERNAL_15;
N_423 <= CPI_DBG_DATA_INTERNAL_16;
N_424 <= CPI_DBG_DATA_INTERNAL_17;
N_425 <= CPI_DBG_DATA_INTERNAL_18;
N_426 <= CPI_DBG_DATA_INTERNAL_19;
N_427 <= CPI_DBG_DATA_INTERNAL_20;
N_428 <= CPI_DBG_DATA_INTERNAL_21;
N_429 <= CPI_DBG_DATA_INTERNAL_22;
N_430 <= CPI_DBG_DATA_INTERNAL_23;
N_431 <= CPI_DBG_DATA_INTERNAL_24;
N_432 <= CPI_DBG_DATA_INTERNAL_25;
N_433 <= CPI_DBG_DATA_INTERNAL_26;
N_434 <= CPI_DBG_DATA_INTERNAL_27;
N_435 <= CPI_DBG_DATA_INTERNAL_28;
N_436 <= CPI_DBG_DATA_INTERNAL_29;
N_437 <= CPI_DBG_DATA_INTERNAL_30;
N_0 <= CPO_DATAZ(0);
N_1_75 <= CPO_DATAZ(1);
N_2_0 <= CPO_DATAZ(2);
N_3_0 <= CPO_DATAZ(3);
N_4_0 <= CPO_DATAZ(4);
N_5_0 <= CPO_DATAZ(5);
N_6_0 <= CPO_DATAZ(6);
N_7_0 <= CPO_DATAZ(7);
N_8_0 <= CPO_DATAZ(8);
N_9_0 <= CPO_DATAZ(9);
N_10_0 <= CPO_DATAZ(10);
N_11_0 <= CPO_DATAZ(11);
N_12_0 <= CPO_DATAZ(12);
N_13_0 <= CPO_DATAZ(13);
N_14_0 <= CPO_DATAZ(14);
N_15_0 <= CPO_DATAZ(15);
N_16_0 <= CPO_DATAZ(16);
N_17_0 <= CPO_DATAZ(17);
N_18_0 <= CPO_DATAZ(18);
N_19_0 <= CPO_DATAZ(19);
N_20_0 <= CPO_DATAZ(20);
N_21_0 <= CPO_DATAZ(21);
N_22_0 <= CPO_DATAZ(22);
N_23_0 <= CPO_DATAZ(23);
N_24_0 <= CPO_DATAZ(24);
N_25_0 <= CPO_DATAZ(25);
N_26_0 <= CPO_DATAZ(26);
N_27_0 <= CPO_DATAZ(27);
N_28_0 <= CPO_DATAZ(28);
N_29_0 <= CPO_DATAZ(29);
N_30_0 <= CPO_DATAZ(30);
N_31_0 <= CPO_DATAZ(31);
N_32_0 <= CPO_EXCZ;
N_33_0 <= CPO_CCZ(0);
N_34_0 <= CPO_CCZ(1);
N_35_0 <= CPO_CCVZ;
N_36_0 <= CPO_LDLOCKZ;
N_37_0 <= CPO_HOLDNZ;
N_38_0 <= CPO_DBG_DATAZ(0);
N_39_0 <= CPO_DBG_DATAZ(1);
N_40_0 <= CPO_DBG_DATAZ(2);
N_41_0 <= CPO_DBG_DATAZ(3);
N_42_0 <= CPO_DBG_DATAZ(4);
N_43_0 <= CPO_DBG_DATAZ(5);
N_44_0 <= CPO_DBG_DATAZ(6);
N_45_0 <= CPO_DBG_DATAZ(7);
N_46_0 <= CPO_DBG_DATAZ(8);
N_47_0 <= CPO_DBG_DATAZ(9);
N_48_0 <= CPO_DBG_DATAZ(10);
N_49_0 <= CPO_DBG_DATAZ(11);
N_50_0 <= CPO_DBG_DATAZ(12);
N_51_0 <= CPO_DBG_DATAZ(13);
N_52_0 <= CPO_DBG_DATAZ(14);
N_53_0 <= CPO_DBG_DATAZ(15);
N_54_0 <= CPO_DBG_DATAZ(16);
N_55_0 <= CPO_DBG_DATAZ(17);
N_56_0 <= CPO_DBG_DATAZ(18);
N_57_0 <= CPO_DBG_DATAZ(19);
N_58_0 <= CPO_DBG_DATAZ(20);
N_59_0 <= CPO_DBG_DATAZ(21);
N_60_0 <= CPO_DBG_DATAZ(22);
N_61_0 <= CPO_DBG_DATAZ(23);
N_62_0 <= CPO_DBG_DATAZ(24);
N_63_0 <= CPO_DBG_DATAZ(25);
N_64_0 <= CPO_DBG_DATAZ(26);
N_65_0 <= CPO_DBG_DATAZ(27);
N_66_0 <= CPO_DBG_DATAZ(28);
N_67_0 <= CPO_DBG_DATAZ(29);
N_68_0 <= CPO_DBG_DATAZ(30);
N_69_0 <= CPO_DBG_DATAZ(31);
N_70_0 <= RFI2_RD1ADDRZ(0);
N_71_0 <= RFI2_RD1ADDRZ(1);
N_72_0 <= RFI2_RD1ADDRZ(2);
N_73_0 <= RFI2_RD1ADDRZ(3);
N_74_0 <= RFI2_RD2ADDRZ(0);
N_75_0 <= RFI2_RD2ADDRZ(1);
N_76_0 <= RFI2_RD2ADDRZ(2);
N_77_0 <= RFI2_RD2ADDRZ(3);
N_78_0 <= RFI2_WRADDRZ(0);
N_79_0 <= RFI2_WRADDRZ(1);
N_80_0 <= RFI2_WRADDRZ(2);
N_81_0 <= RFI2_WRADDRZ(3);
N_82_0 <= RFI1_WRDATAZ(0);
N_83_0 <= RFI1_WRDATAZ(1);
N_84_0 <= RFI1_WRDATAZ(2);
N_85_0 <= RFI1_WRDATAZ(3);
N_86_0 <= RFI1_WRDATAZ(4);
N_87_0 <= RFI1_WRDATAZ(5);
N_88_0 <= RFI1_WRDATAZ(6);
N_89_0 <= RFI1_WRDATAZ(7);
N_90_0 <= RFI1_WRDATAZ(8);
N_91_0 <= RFI1_WRDATAZ(9);
N_92_0 <= RFI1_WRDATAZ(10);
N_93_0 <= RFI1_WRDATAZ(11);
N_94_0 <= RFI1_WRDATAZ(12);
N_95_0 <= RFI1_WRDATAZ(13);
N_96_0 <= RFI1_WRDATAZ(14);
N_97_0 <= RFI1_WRDATAZ(15);
N_98_0 <= RFI1_WRDATAZ(16);
N_99_0 <= RFI1_WRDATAZ(17);
N_100_0 <= RFI1_WRDATAZ(18);
N_101_0 <= RFI1_WRDATAZ(19);
N_102_0 <= RFI1_WRDATAZ(20);
N_103_0 <= RFI1_WRDATAZ(21);
N_104_0 <= RFI1_WRDATAZ(22);
N_105_0 <= RFI1_WRDATAZ(23);
N_106_0 <= RFI1_WRDATAZ(24);
N_107_0 <= RFI1_WRDATAZ(25);
N_108_0 <= RFI1_WRDATAZ(26);
N_109_0 <= RFI1_WRDATAZ(27);
N_110_0 <= RFI1_WRDATAZ(28);
N_111_0 <= RFI1_WRDATAZ(29);
N_112_0 <= RFI1_WRDATAZ(30);
N_113_0 <= RFI1_WRDATAZ(31);
N_114_0 <= RFI1_REN1Z;
N_115_0 <= RFI1_REN2Z;
N_116_0 <= RFI1_WRENZ;
N_117_0 <= RFI2_RD1ADDRZ(0);
N_118_0 <= RFI2_RD1ADDRZ(1);
N_119_0 <= RFI2_RD1ADDRZ(2);
N_120_0 <= RFI2_RD1ADDRZ(3);
N_121_0 <= RFI2_RD2ADDRZ(0);
N_122_0 <= RFI2_RD2ADDRZ(1);
N_123_0 <= RFI2_RD2ADDRZ(2);
N_124_0 <= RFI2_RD2ADDRZ(3);
N_125_0 <= RFI2_WRADDRZ(0);
N_126_0 <= RFI2_WRADDRZ(1);
N_127_0 <= RFI2_WRADDRZ(2);
N_128_0 <= RFI2_WRADDRZ(3);
N_129_0 <= RFI2_WRDATAZ(0);
N_130_0 <= RFI2_WRDATAZ(1);
N_131_0 <= RFI2_WRDATAZ(2);
N_132_0 <= RFI2_WRDATAZ(3);
N_133_0 <= RFI2_WRDATAZ(4);
N_134_0 <= RFI2_WRDATAZ(5);
N_135_0 <= RFI2_WRDATAZ(6);
N_136_0 <= RFI2_WRDATAZ(7);
N_137_0 <= RFI2_WRDATAZ(8);
N_138_0 <= RFI2_WRDATAZ(9);
N_139_0 <= RFI2_WRDATAZ(10);
N_140_0 <= RFI2_WRDATAZ(11);
N_141_0 <= RFI2_WRDATAZ(12);
N_142_0 <= RFI2_WRDATAZ(13);
N_143_0 <= RFI2_WRDATAZ(14);
N_144_0 <= RFI2_WRDATAZ(15);
N_145_0 <= RFI2_WRDATAZ(16);
N_146_0 <= RFI2_WRDATAZ(17);
N_147_0 <= RFI2_WRDATAZ(18);
N_148_0 <= RFI2_WRDATAZ(19);
N_149_0 <= RFI2_WRDATAZ(20);
N_150_0 <= RFI2_WRDATAZ(21);
N_151_0 <= RFI2_WRDATAZ(22);
N_152_0 <= RFI2_WRDATAZ(23);
N_153_0 <= RFI2_WRDATAZ(24);
N_154_0 <= RFI2_WRDATAZ(25);
N_155_0 <= RFI2_WRDATAZ(26);
N_156_0 <= RFI2_WRDATAZ(27);
N_157_0 <= RFI2_WRDATAZ(28);
N_158_0 <= RFI2_WRDATAZ(29);
N_159_0 <= RFI2_WRDATAZ(30);
N_160_0 <= RFI2_WRDATAZ(31);
N_161_0 <= RFI2_REN1Z;
N_162_0 <= RFI2_REN2Z;
N_163_0 <= RFI2_WRENZ;
N_602 <= RFO1_DATA1_INTERNAL;
N_603 <= RFO1_DATA1_INTERNAL_0;
N_604 <= RFO1_DATA1_INTERNAL_1;
N_605 <= RFO1_DATA1_INTERNAL_2;
N_606 <= RFO1_DATA1_INTERNAL_3;
N_607 <= RFO1_DATA1_INTERNAL_4;
N_608 <= RFO1_DATA1_INTERNAL_5;
N_609 <= RFO1_DATA1_INTERNAL_6;
N_610 <= RFO1_DATA1_INTERNAL_7;
N_611 <= RFO1_DATA1_INTERNAL_8;
N_612 <= RFO1_DATA1_INTERNAL_9;
N_613 <= RFO1_DATA1_INTERNAL_10;
N_614 <= RFO1_DATA1_INTERNAL_11;
N_615 <= RFO1_DATA1_INTERNAL_12;
N_616 <= RFO1_DATA1_INTERNAL_13;
N_617 <= RFO1_DATA1_INTERNAL_14;
N_618 <= RFO1_DATA1_INTERNAL_15;
N_619 <= RFO1_DATA1_INTERNAL_16;
N_620 <= RFO1_DATA1_INTERNAL_17;
N_621 <= RFO1_DATA1_INTERNAL_18;
N_622 <= RFO1_DATA1_INTERNAL_19;
N_623 <= RFO1_DATA1_INTERNAL_20;
N_624 <= RFO1_DATA1_INTERNAL_21;
N_625 <= RFO1_DATA1_INTERNAL_22;
N_626 <= RFO1_DATA1_INTERNAL_23;
N_627 <= RFO1_DATA1_INTERNAL_24;
N_628 <= RFO1_DATA1_INTERNAL_25;
N_629 <= RFO1_DATA1_INTERNAL_26;
N_630 <= RFO1_DATA1_INTERNAL_27;
N_631 <= RFO1_DATA1_INTERNAL_28;
N_632 <= RFO1_DATA1_INTERNAL_29;
N_633 <= RFO1_DATA1_INTERNAL_30;
N_634 <= RFO1_DATA2_INTERNAL;
N_635 <= RFO1_DATA2_INTERNAL_0;
N_636 <= RFO1_DATA2_INTERNAL_1;
N_637 <= RFO1_DATA2_INTERNAL_2;
N_638 <= RFO1_DATA2_INTERNAL_3;
N_639 <= RFO1_DATA2_INTERNAL_4;
N_640 <= RFO1_DATA2_INTERNAL_5;
N_641 <= RFO1_DATA2_INTERNAL_6;
N_642 <= RFO1_DATA2_INTERNAL_7;
N_643 <= RFO1_DATA2_INTERNAL_8;
N_644 <= RFO1_DATA2_INTERNAL_9;
N_645 <= RFO1_DATA2_INTERNAL_10;
N_646 <= RFO1_DATA2_INTERNAL_11;
N_647 <= RFO1_DATA2_INTERNAL_12;
N_648 <= RFO1_DATA2_INTERNAL_13;
N_649 <= RFO1_DATA2_INTERNAL_14;
N_650 <= RFO1_DATA2_INTERNAL_15;
N_651 <= RFO1_DATA2_INTERNAL_16;
N_652 <= RFO1_DATA2_INTERNAL_17;
N_653 <= RFO1_DATA2_INTERNAL_18;
N_654 <= RFO1_DATA2_INTERNAL_19;
N_655 <= RFO1_DATA2_INTERNAL_20;
N_656 <= RFO1_DATA2_INTERNAL_21;
N_657 <= RFO1_DATA2_INTERNAL_22;
N_658 <= RFO1_DATA2_INTERNAL_23;
N_659 <= RFO1_DATA2_INTERNAL_24;
N_660 <= RFO1_DATA2_INTERNAL_25;
N_661 <= RFO1_DATA2_INTERNAL_26;
N_662 <= RFO1_DATA2_INTERNAL_27;
N_663 <= RFO1_DATA2_INTERNAL_28;
N_664 <= RFO1_DATA2_INTERNAL_29;
N_665 <= RFO1_DATA2_INTERNAL_30;
N_666 <= RFO2_DATA1_INTERNAL;
N_667 <= RFO2_DATA1_INTERNAL_0;
N_668 <= RFO2_DATA1_INTERNAL_1;
N_669 <= RFO2_DATA1_INTERNAL_2;
N_670 <= RFO2_DATA1_INTERNAL_3;
N_671 <= RFO2_DATA1_INTERNAL_4;
N_672 <= RFO2_DATA1_INTERNAL_5;
N_673 <= RFO2_DATA1_INTERNAL_6;
N_674 <= RFO2_DATA1_INTERNAL_7;
N_675 <= RFO2_DATA1_INTERNAL_8;
N_676 <= RFO2_DATA1_INTERNAL_9;
N_677 <= RFO2_DATA1_INTERNAL_10;
N_678 <= RFO2_DATA1_INTERNAL_11;
N_679 <= RFO2_DATA1_INTERNAL_12;
N_680 <= RFO2_DATA1_INTERNAL_13;
N_681 <= RFO2_DATA1_INTERNAL_14;
N_682 <= RFO2_DATA1_INTERNAL_15;
N_683 <= RFO2_DATA1_INTERNAL_16;
N_684 <= RFO2_DATA1_INTERNAL_17;
N_685 <= RFO2_DATA1_INTERNAL_18;
N_686 <= RFO2_DATA1_INTERNAL_19;
N_687 <= RFO2_DATA1_INTERNAL_20;
N_688 <= RFO2_DATA1_INTERNAL_21;
N_689 <= RFO2_DATA1_INTERNAL_22;
N_690 <= RFO2_DATA1_INTERNAL_23;
N_691 <= RFO2_DATA1_INTERNAL_24;
N_692 <= RFO2_DATA1_INTERNAL_25;
N_693 <= RFO2_DATA1_INTERNAL_26;
N_694 <= RFO2_DATA1_INTERNAL_27;
N_695 <= RFO2_DATA1_INTERNAL_28;
N_696 <= RFO2_DATA1_INTERNAL_29;
N_697 <= RFO2_DATA1_INTERNAL_30;
N_698 <= RFO2_DATA2_INTERNAL;
N_699 <= RFO2_DATA2_INTERNAL_0;
N_700 <= RFO2_DATA2_INTERNAL_1;
N_701 <= RFO2_DATA2_INTERNAL_2;
N_702 <= RFO2_DATA2_INTERNAL_3;
N_703 <= RFO2_DATA2_INTERNAL_4;
N_704 <= RFO2_DATA2_INTERNAL_5;
N_705 <= RFO2_DATA2_INTERNAL_6;
N_706 <= RFO2_DATA2_INTERNAL_7;
N_707 <= RFO2_DATA2_INTERNAL_8;
N_708 <= RFO2_DATA2_INTERNAL_9;
N_709 <= RFO2_DATA2_INTERNAL_10;
N_710 <= RFO2_DATA2_INTERNAL_11;
N_711 <= RFO2_DATA2_INTERNAL_12;
N_712 <= RFO2_DATA2_INTERNAL_13;
N_713 <= RFO2_DATA2_INTERNAL_14;
N_714 <= RFO2_DATA2_INTERNAL_15;
N_715 <= RFO2_DATA2_INTERNAL_16;
N_716 <= RFO2_DATA2_INTERNAL_17;
N_717 <= RFO2_DATA2_INTERNAL_18;
N_718 <= RFO2_DATA2_INTERNAL_19;
N_719 <= RFO2_DATA2_INTERNAL_20;
N_720 <= RFO2_DATA2_INTERNAL_21;
N_721 <= RFO2_DATA2_INTERNAL_22;
N_722 <= RFO2_DATA2_INTERNAL_23;
N_723 <= RFO2_DATA2_INTERNAL_24;
N_724 <= RFO2_DATA2_INTERNAL_25;
N_725 <= RFO2_DATA2_INTERNAL_26;
N_726 <= RFO2_DATA2_INTERNAL_27;
N_727 <= RFO2_DATA2_INTERNAL_28;
N_728 <= RFO2_DATA2_INTERNAL_29;
N_729 <= RFO2_DATA2_INTERNAL_30;
cpo_data(0) <= N_0;
cpo_data(1) <= N_1_75;
cpo_data(2) <= N_2_0;
cpo_data(3) <= N_3_0;
cpo_data(4) <= N_4_0;
cpo_data(5) <= N_5_0;
cpo_data(6) <= N_6_0;
cpo_data(7) <= N_7_0;
cpo_data(8) <= N_8_0;
cpo_data(9) <= N_9_0;
cpo_data(10) <= N_10_0;
cpo_data(11) <= N_11_0;
cpo_data(12) <= N_12_0;
cpo_data(13) <= N_13_0;
cpo_data(14) <= N_14_0;
cpo_data(15) <= N_15_0;
cpo_data(16) <= N_16_0;
cpo_data(17) <= N_17_0;
cpo_data(18) <= N_18_0;
cpo_data(19) <= N_19_0;
cpo_data(20) <= N_20_0;
cpo_data(21) <= N_21_0;
cpo_data(22) <= N_22_0;
cpo_data(23) <= N_23_0;
cpo_data(24) <= N_24_0;
cpo_data(25) <= N_25_0;
cpo_data(26) <= N_26_0;
cpo_data(27) <= N_27_0;
cpo_data(28) <= N_28_0;
cpo_data(29) <= N_29_0;
cpo_data(30) <= N_30_0;
cpo_data(31) <= N_31_0;
cpo_exc <= N_32_0;
cpo_cc(0) <= N_33_0;
cpo_cc(1) <= N_34_0;
cpo_ccv <= N_35_0;
cpo_ldlock <= N_36_0;
cpo_holdn <= N_37_0;
cpo_dbg_data(0) <= N_38_0;
cpo_dbg_data(1) <= N_39_0;
cpo_dbg_data(2) <= N_40_0;
cpo_dbg_data(3) <= N_41_0;
cpo_dbg_data(4) <= N_42_0;
cpo_dbg_data(5) <= N_43_0;
cpo_dbg_data(6) <= N_44_0;
cpo_dbg_data(7) <= N_45_0;
cpo_dbg_data(8) <= N_46_0;
cpo_dbg_data(9) <= N_47_0;
cpo_dbg_data(10) <= N_48_0;
cpo_dbg_data(11) <= N_49_0;
cpo_dbg_data(12) <= N_50_0;
cpo_dbg_data(13) <= N_51_0;
cpo_dbg_data(14) <= N_52_0;
cpo_dbg_data(15) <= N_53_0;
cpo_dbg_data(16) <= N_54_0;
cpo_dbg_data(17) <= N_55_0;
cpo_dbg_data(18) <= N_56_0;
cpo_dbg_data(19) <= N_57_0;
cpo_dbg_data(20) <= N_58_0;
cpo_dbg_data(21) <= N_59_0;
cpo_dbg_data(22) <= N_60_0;
cpo_dbg_data(23) <= N_61_0;
cpo_dbg_data(24) <= N_62_0;
cpo_dbg_data(25) <= N_63_0;
cpo_dbg_data(26) <= N_64_0;
cpo_dbg_data(27) <= N_65_0;
cpo_dbg_data(28) <= N_66_0;
cpo_dbg_data(29) <= N_67_0;
cpo_dbg_data(30) <= N_68_0;
cpo_dbg_data(31) <= N_69_0;
rfi1_rd1addr(0) <= N_70_0;
rfi1_rd1addr(1) <= N_71_0;
rfi1_rd1addr(2) <= N_72_0;
rfi1_rd1addr(3) <= N_73_0;
rfi1_rd2addr(0) <= N_74_0;
rfi1_rd2addr(1) <= N_75_0;
rfi1_rd2addr(2) <= N_76_0;
rfi1_rd2addr(3) <= N_77_0;
rfi1_wraddr(0) <= N_78_0;
rfi1_wraddr(1) <= N_79_0;
rfi1_wraddr(2) <= N_80_0;
rfi1_wraddr(3) <= N_81_0;
rfi1_wrdata(0) <= N_82_0;
rfi1_wrdata(1) <= N_83_0;
rfi1_wrdata(2) <= N_84_0;
rfi1_wrdata(3) <= N_85_0;
rfi1_wrdata(4) <= N_86_0;
rfi1_wrdata(5) <= N_87_0;
rfi1_wrdata(6) <= N_88_0;
rfi1_wrdata(7) <= N_89_0;
rfi1_wrdata(8) <= N_90_0;
rfi1_wrdata(9) <= N_91_0;
rfi1_wrdata(10) <= N_92_0;
rfi1_wrdata(11) <= N_93_0;
rfi1_wrdata(12) <= N_94_0;
rfi1_wrdata(13) <= N_95_0;
rfi1_wrdata(14) <= N_96_0;
rfi1_wrdata(15) <= N_97_0;
rfi1_wrdata(16) <= N_98_0;
rfi1_wrdata(17) <= N_99_0;
rfi1_wrdata(18) <= N_100_0;
rfi1_wrdata(19) <= N_101_0;
rfi1_wrdata(20) <= N_102_0;
rfi1_wrdata(21) <= N_103_0;
rfi1_wrdata(22) <= N_104_0;
rfi1_wrdata(23) <= N_105_0;
rfi1_wrdata(24) <= N_106_0;
rfi1_wrdata(25) <= N_107_0;
rfi1_wrdata(26) <= N_108_0;
rfi1_wrdata(27) <= N_109_0;
rfi1_wrdata(28) <= N_110_0;
rfi1_wrdata(29) <= N_111_0;
rfi1_wrdata(30) <= N_112_0;
rfi1_wrdata(31) <= N_113_0;
rfi1_ren1 <= N_114_0;
rfi1_ren2 <= N_115_0;
rfi1_wren <= N_116_0;
rfi2_rd1addr(0) <= N_117_0;
rfi2_rd1addr(1) <= N_118_0;
rfi2_rd1addr(2) <= N_119_0;
rfi2_rd1addr(3) <= N_120_0;
rfi2_rd2addr(0) <= N_121_0;
rfi2_rd2addr(1) <= N_122_0;
rfi2_rd2addr(2) <= N_123_0;
rfi2_rd2addr(3) <= N_124_0;
rfi2_wraddr(0) <= N_125_0;
rfi2_wraddr(1) <= N_126_0;
rfi2_wraddr(2) <= N_127_0;
rfi2_wraddr(3) <= N_128_0;
rfi2_wrdata(0) <= N_129_0;
rfi2_wrdata(1) <= N_130_0;
rfi2_wrdata(2) <= N_131_0;
rfi2_wrdata(3) <= N_132_0;
rfi2_wrdata(4) <= N_133_0;
rfi2_wrdata(5) <= N_134_0;
rfi2_wrdata(6) <= N_135_0;
rfi2_wrdata(7) <= N_136_0;
rfi2_wrdata(8) <= N_137_0;
rfi2_wrdata(9) <= N_138_0;
rfi2_wrdata(10) <= N_139_0;
rfi2_wrdata(11) <= N_140_0;
rfi2_wrdata(12) <= N_141_0;
rfi2_wrdata(13) <= N_142_0;
rfi2_wrdata(14) <= N_143_0;
rfi2_wrdata(15) <= N_144_0;
rfi2_wrdata(16) <= N_145_0;
rfi2_wrdata(17) <= N_146_0;
rfi2_wrdata(18) <= N_147_0;
rfi2_wrdata(19) <= N_148_0;
rfi2_wrdata(20) <= N_149_0;
rfi2_wrdata(21) <= N_150_0;
rfi2_wrdata(22) <= N_151_0;
rfi2_wrdata(23) <= N_152_0;
rfi2_wrdata(24) <= N_153_0;
rfi2_wrdata(25) <= N_154_0;
rfi2_wrdata(26) <= N_155_0;
rfi2_wrdata(27) <= N_156_0;
rfi2_wrdata(28) <= N_157_0;
rfi2_wrdata(29) <= N_158_0;
rfi2_wrdata(30) <= N_159_0;
rfi2_wrdata(31) <= N_160_0;
rfi2_ren1 <= N_161_0;
rfi2_ren2 <= N_162_0;
rfi2_wren <= N_163_0;
RST_INTERNAL <= rst;
CLK_INTERNAL <= clk;
HOLDN_INTERNAL <= holdn;
CPI_FLUSH_INTERNAL <= cpi_flush;
CPI_EXACK_INTERNAL <= cpi_exack;
CPI_A_RS1_INTERNAL <= cpi_a_rs1(0);
CPI_A_RS1_INTERNAL_0 <= cpi_a_rs1(1);
CPI_A_RS1_INTERNAL_1 <= cpi_a_rs1(2);
CPI_A_RS1_INTERNAL_2 <= cpi_a_rs1(3);
CPI_A_RS1_INTERNAL_3 <= cpi_a_rs1(4);
CPI_D_PC_INTERNAL <= cpi_d_pc(0);
CPI_D_PC_INTERNAL_0 <= cpi_d_pc(1);
CPI_D_PC_INTERNAL_1 <= cpi_d_pc(2);
CPI_D_PC_INTERNAL_2 <= cpi_d_pc(3);
CPI_D_PC_INTERNAL_3 <= cpi_d_pc(4);
CPI_D_PC_INTERNAL_4 <= cpi_d_pc(5);
CPI_D_PC_INTERNAL_5 <= cpi_d_pc(6);
CPI_D_PC_INTERNAL_6 <= cpi_d_pc(7);
CPI_D_PC_INTERNAL_7 <= cpi_d_pc(8);
CPI_D_PC_INTERNAL_8 <= cpi_d_pc(9);
CPI_D_PC_INTERNAL_9 <= cpi_d_pc(10);
CPI_D_PC_INTERNAL_10 <= cpi_d_pc(11);
CPI_D_PC_INTERNAL_11 <= cpi_d_pc(12);
CPI_D_PC_INTERNAL_12 <= cpi_d_pc(13);
CPI_D_PC_INTERNAL_13 <= cpi_d_pc(14);
CPI_D_PC_INTERNAL_14 <= cpi_d_pc(15);
CPI_D_PC_INTERNAL_15 <= cpi_d_pc(16);
CPI_D_PC_INTERNAL_16 <= cpi_d_pc(17);
CPI_D_PC_INTERNAL_17 <= cpi_d_pc(18);
CPI_D_PC_INTERNAL_18 <= cpi_d_pc(19);
CPI_D_PC_INTERNAL_19 <= cpi_d_pc(20);
CPI_D_PC_INTERNAL_20 <= cpi_d_pc(21);
CPI_D_PC_INTERNAL_21 <= cpi_d_pc(22);
CPI_D_PC_INTERNAL_22 <= cpi_d_pc(23);
CPI_D_PC_INTERNAL_23 <= cpi_d_pc(24);
CPI_D_PC_INTERNAL_24 <= cpi_d_pc(25);
CPI_D_PC_INTERNAL_25 <= cpi_d_pc(26);
CPI_D_PC_INTERNAL_26 <= cpi_d_pc(27);
CPI_D_PC_INTERNAL_27 <= cpi_d_pc(28);
CPI_D_PC_INTERNAL_28 <= cpi_d_pc(29);
CPI_D_PC_INTERNAL_29 <= cpi_d_pc(30);
CPI_D_PC_INTERNAL_30 <= cpi_d_pc(31);
CPI_D_INST_INTERNAL <= cpi_d_inst(0);
CPI_D_INST_INTERNAL_0 <= cpi_d_inst(1);
CPI_D_INST_INTERNAL_1 <= cpi_d_inst(2);
CPI_D_INST_INTERNAL_2 <= cpi_d_inst(3);
CPI_D_INST_INTERNAL_3 <= cpi_d_inst(4);
CPI_D_INST_INTERNAL_4 <= cpi_d_inst(5);
CPI_D_INST_INTERNAL_5 <= cpi_d_inst(6);
CPI_D_INST_INTERNAL_6 <= cpi_d_inst(7);
CPI_D_INST_INTERNAL_7 <= cpi_d_inst(8);
CPI_D_INST_INTERNAL_8 <= cpi_d_inst(9);
CPI_D_INST_INTERNAL_9 <= cpi_d_inst(10);
CPI_D_INST_INTERNAL_10 <= cpi_d_inst(11);
CPI_D_INST_INTERNAL_11 <= cpi_d_inst(12);
CPI_D_INST_INTERNAL_12 <= cpi_d_inst(13);
CPI_D_INST_INTERNAL_13 <= cpi_d_inst(14);
CPI_D_INST_INTERNAL_14 <= cpi_d_inst(15);
CPI_D_INST_INTERNAL_15 <= cpi_d_inst(16);
CPI_D_INST_INTERNAL_16 <= cpi_d_inst(17);
CPI_D_INST_INTERNAL_17 <= cpi_d_inst(18);
CPI_D_INST_INTERNAL_18 <= cpi_d_inst(19);
CPI_D_INST_INTERNAL_19 <= cpi_d_inst(20);
CPI_D_INST_INTERNAL_20 <= cpi_d_inst(21);
CPI_D_INST_INTERNAL_21 <= cpi_d_inst(22);
CPI_D_INST_INTERNAL_22 <= cpi_d_inst(23);
CPI_D_INST_INTERNAL_23 <= cpi_d_inst(24);
CPI_D_INST_INTERNAL_24 <= cpi_d_inst(25);
CPI_D_INST_INTERNAL_25 <= cpi_d_inst(26);
CPI_D_INST_INTERNAL_26 <= cpi_d_inst(27);
CPI_D_INST_INTERNAL_27 <= cpi_d_inst(28);
CPI_D_INST_INTERNAL_28 <= cpi_d_inst(29);
CPI_D_INST_INTERNAL_29 <= cpi_d_inst(30);
CPI_D_INST_INTERNAL_30 <= cpi_d_inst(31);
CPI_D_CNT_INTERNAL <= cpi_d_cnt(0);
CPI_D_CNT_INTERNAL_0 <= cpi_d_cnt(1);
CPI_D_TRAP_INTERNAL <= cpi_d_trap;
CPI_D_ANNUL_INTERNAL <= cpi_d_annul;
CPI_D_PV_INTERNAL <= cpi_d_pv;
CPI_A_PC_INTERNAL <= cpi_a_pc(0);
CPI_A_PC_INTERNAL_0 <= cpi_a_pc(1);
CPI_A_PC_INTERNAL_1 <= cpi_a_pc(2);
CPI_A_PC_INTERNAL_2 <= cpi_a_pc(3);
CPI_A_PC_INTERNAL_3 <= cpi_a_pc(4);
CPI_A_PC_INTERNAL_4 <= cpi_a_pc(5);
CPI_A_PC_INTERNAL_5 <= cpi_a_pc(6);
CPI_A_PC_INTERNAL_6 <= cpi_a_pc(7);
CPI_A_PC_INTERNAL_7 <= cpi_a_pc(8);
CPI_A_PC_INTERNAL_8 <= cpi_a_pc(9);
CPI_A_PC_INTERNAL_9 <= cpi_a_pc(10);
CPI_A_PC_INTERNAL_10 <= cpi_a_pc(11);
CPI_A_PC_INTERNAL_11 <= cpi_a_pc(12);
CPI_A_PC_INTERNAL_12 <= cpi_a_pc(13);
CPI_A_PC_INTERNAL_13 <= cpi_a_pc(14);
CPI_A_PC_INTERNAL_14 <= cpi_a_pc(15);
CPI_A_PC_INTERNAL_15 <= cpi_a_pc(16);
CPI_A_PC_INTERNAL_16 <= cpi_a_pc(17);
CPI_A_PC_INTERNAL_17 <= cpi_a_pc(18);
CPI_A_PC_INTERNAL_18 <= cpi_a_pc(19);
CPI_A_PC_INTERNAL_19 <= cpi_a_pc(20);
CPI_A_PC_INTERNAL_20 <= cpi_a_pc(21);
CPI_A_PC_INTERNAL_21 <= cpi_a_pc(22);
CPI_A_PC_INTERNAL_22 <= cpi_a_pc(23);
CPI_A_PC_INTERNAL_23 <= cpi_a_pc(24);
CPI_A_PC_INTERNAL_24 <= cpi_a_pc(25);
CPI_A_PC_INTERNAL_25 <= cpi_a_pc(26);
CPI_A_PC_INTERNAL_26 <= cpi_a_pc(27);
CPI_A_PC_INTERNAL_27 <= cpi_a_pc(28);
CPI_A_PC_INTERNAL_28 <= cpi_a_pc(29);
CPI_A_PC_INTERNAL_29 <= cpi_a_pc(30);
CPI_A_PC_INTERNAL_30 <= cpi_a_pc(31);
CPI_A_INST_INTERNAL <= cpi_a_inst(0);
CPI_A_INST_INTERNAL_0 <= cpi_a_inst(1);
CPI_A_INST_INTERNAL_1 <= cpi_a_inst(2);
CPI_A_INST_INTERNAL_2 <= cpi_a_inst(3);
CPI_A_INST_INTERNAL_3 <= cpi_a_inst(4);
CPI_A_INST_INTERNAL_4 <= cpi_a_inst(5);
CPI_A_INST_INTERNAL_5 <= cpi_a_inst(6);
CPI_A_INST_INTERNAL_6 <= cpi_a_inst(7);
CPI_A_INST_INTERNAL_7 <= cpi_a_inst(8);
CPI_A_INST_INTERNAL_8 <= cpi_a_inst(9);
CPI_A_INST_INTERNAL_9 <= cpi_a_inst(10);
CPI_A_INST_INTERNAL_10 <= cpi_a_inst(11);
CPI_A_INST_INTERNAL_11 <= cpi_a_inst(12);
CPI_A_INST_INTERNAL_12 <= cpi_a_inst(13);
CPI_A_INST_INTERNAL_13 <= cpi_a_inst(14);
CPI_A_INST_INTERNAL_14 <= cpi_a_inst(15);
CPI_A_INST_INTERNAL_15 <= cpi_a_inst(16);
CPI_A_INST_INTERNAL_16 <= cpi_a_inst(17);
CPI_A_INST_INTERNAL_17 <= cpi_a_inst(18);
CPI_A_INST_INTERNAL_18 <= cpi_a_inst(19);
CPI_A_INST_INTERNAL_19 <= cpi_a_inst(20);
CPI_A_INST_INTERNAL_20 <= cpi_a_inst(21);
CPI_A_INST_INTERNAL_21 <= cpi_a_inst(22);
CPI_A_INST_INTERNAL_22 <= cpi_a_inst(23);
CPI_A_INST_INTERNAL_23 <= cpi_a_inst(24);
CPI_A_INST_INTERNAL_24 <= cpi_a_inst(25);
CPI_A_INST_INTERNAL_25 <= cpi_a_inst(26);
CPI_A_INST_INTERNAL_26 <= cpi_a_inst(27);
CPI_A_INST_INTERNAL_27 <= cpi_a_inst(28);
CPI_A_INST_INTERNAL_28 <= cpi_a_inst(29);
CPI_A_INST_INTERNAL_29 <= cpi_a_inst(30);
CPI_A_INST_INTERNAL_30 <= cpi_a_inst(31);
CPI_A_CNT_INTERNAL <= cpi_a_cnt(0);
CPI_A_CNT_INTERNAL_0 <= cpi_a_cnt(1);
CPI_A_TRAP_INTERNAL <= cpi_a_trap;
CPI_A_ANNUL_INTERNAL <= cpi_a_annul;
CPI_A_PV_INTERNAL <= cpi_a_pv;
CPI_E_PC_INTERNAL <= cpi_e_pc(0);
CPI_E_PC_INTERNAL_0 <= cpi_e_pc(1);
CPI_E_PC_INTERNAL_1 <= cpi_e_pc(2);
CPI_E_PC_INTERNAL_2 <= cpi_e_pc(3);
CPI_E_PC_INTERNAL_3 <= cpi_e_pc(4);
CPI_E_PC_INTERNAL_4 <= cpi_e_pc(5);
CPI_E_PC_INTERNAL_5 <= cpi_e_pc(6);
CPI_E_PC_INTERNAL_6 <= cpi_e_pc(7);
CPI_E_PC_INTERNAL_7 <= cpi_e_pc(8);
CPI_E_PC_INTERNAL_8 <= cpi_e_pc(9);
CPI_E_PC_INTERNAL_9 <= cpi_e_pc(10);
CPI_E_PC_INTERNAL_10 <= cpi_e_pc(11);
CPI_E_PC_INTERNAL_11 <= cpi_e_pc(12);
CPI_E_PC_INTERNAL_12 <= cpi_e_pc(13);
CPI_E_PC_INTERNAL_13 <= cpi_e_pc(14);
CPI_E_PC_INTERNAL_14 <= cpi_e_pc(15);
CPI_E_PC_INTERNAL_15 <= cpi_e_pc(16);
CPI_E_PC_INTERNAL_16 <= cpi_e_pc(17);
CPI_E_PC_INTERNAL_17 <= cpi_e_pc(18);
CPI_E_PC_INTERNAL_18 <= cpi_e_pc(19);
CPI_E_PC_INTERNAL_19 <= cpi_e_pc(20);
CPI_E_PC_INTERNAL_20 <= cpi_e_pc(21);
CPI_E_PC_INTERNAL_21 <= cpi_e_pc(22);
CPI_E_PC_INTERNAL_22 <= cpi_e_pc(23);
CPI_E_PC_INTERNAL_23 <= cpi_e_pc(24);
CPI_E_PC_INTERNAL_24 <= cpi_e_pc(25);
CPI_E_PC_INTERNAL_25 <= cpi_e_pc(26);
CPI_E_PC_INTERNAL_26 <= cpi_e_pc(27);
CPI_E_PC_INTERNAL_27 <= cpi_e_pc(28);
CPI_E_PC_INTERNAL_28 <= cpi_e_pc(29);
CPI_E_PC_INTERNAL_29 <= cpi_e_pc(30);
CPI_E_PC_INTERNAL_30 <= cpi_e_pc(31);
CPI_E_INST_INTERNAL <= cpi_e_inst(0);
CPI_E_INST_INTERNAL_0 <= cpi_e_inst(1);
CPI_E_INST_INTERNAL_1 <= cpi_e_inst(2);
CPI_E_INST_INTERNAL_2 <= cpi_e_inst(3);
CPI_E_INST_INTERNAL_3 <= cpi_e_inst(4);
CPI_E_INST_INTERNAL_4 <= cpi_e_inst(5);
CPI_E_INST_INTERNAL_5 <= cpi_e_inst(6);
CPI_E_INST_INTERNAL_6 <= cpi_e_inst(7);
CPI_E_INST_INTERNAL_7 <= cpi_e_inst(8);
CPI_E_INST_INTERNAL_8 <= cpi_e_inst(9);
CPI_E_INST_INTERNAL_9 <= cpi_e_inst(10);
CPI_E_INST_INTERNAL_10 <= cpi_e_inst(11);
CPI_E_INST_INTERNAL_11 <= cpi_e_inst(12);
CPI_E_INST_INTERNAL_12 <= cpi_e_inst(13);
CPI_E_INST_INTERNAL_13 <= cpi_e_inst(14);
CPI_E_INST_INTERNAL_14 <= cpi_e_inst(15);
CPI_E_INST_INTERNAL_15 <= cpi_e_inst(16);
CPI_E_INST_INTERNAL_16 <= cpi_e_inst(17);
CPI_E_INST_INTERNAL_17 <= cpi_e_inst(18);
CPI_E_INST_INTERNAL_18 <= cpi_e_inst(19);
CPI_E_INST_INTERNAL_19 <= cpi_e_inst(20);
CPI_E_INST_INTERNAL_20 <= cpi_e_inst(21);
CPI_E_INST_INTERNAL_21 <= cpi_e_inst(22);
CPI_E_INST_INTERNAL_22 <= cpi_e_inst(23);
CPI_E_INST_INTERNAL_23 <= cpi_e_inst(24);
CPI_E_INST_INTERNAL_24 <= cpi_e_inst(25);
CPI_E_INST_INTERNAL_25 <= cpi_e_inst(26);
CPI_E_INST_INTERNAL_26 <= cpi_e_inst(27);
CPI_E_INST_INTERNAL_27 <= cpi_e_inst(28);
CPI_E_INST_INTERNAL_28 <= cpi_e_inst(29);
CPI_E_INST_INTERNAL_29 <= cpi_e_inst(30);
CPI_E_INST_INTERNAL_30 <= cpi_e_inst(31);
CPI_E_CNT_INTERNAL <= cpi_e_cnt(0);
CPI_E_CNT_INTERNAL_0 <= cpi_e_cnt(1);
CPI_E_TRAP_INTERNAL <= cpi_e_trap;
CPI_E_ANNUL_INTERNAL <= cpi_e_annul;
CPI_E_PV_INTERNAL <= cpi_e_pv;
CPI_M_PC_INTERNAL <= cpi_m_pc(0);
CPI_M_PC_INTERNAL_0 <= cpi_m_pc(1);
CPI_M_PC_INTERNAL_1 <= cpi_m_pc(2);
CPI_M_PC_INTERNAL_2 <= cpi_m_pc(3);
CPI_M_PC_INTERNAL_3 <= cpi_m_pc(4);
CPI_M_PC_INTERNAL_4 <= cpi_m_pc(5);
CPI_M_PC_INTERNAL_5 <= cpi_m_pc(6);
CPI_M_PC_INTERNAL_6 <= cpi_m_pc(7);
CPI_M_PC_INTERNAL_7 <= cpi_m_pc(8);
CPI_M_PC_INTERNAL_8 <= cpi_m_pc(9);
CPI_M_PC_INTERNAL_9 <= cpi_m_pc(10);
CPI_M_PC_INTERNAL_10 <= cpi_m_pc(11);
CPI_M_PC_INTERNAL_11 <= cpi_m_pc(12);
CPI_M_PC_INTERNAL_12 <= cpi_m_pc(13);
CPI_M_PC_INTERNAL_13 <= cpi_m_pc(14);
CPI_M_PC_INTERNAL_14 <= cpi_m_pc(15);
CPI_M_PC_INTERNAL_15 <= cpi_m_pc(16);
CPI_M_PC_INTERNAL_16 <= cpi_m_pc(17);
CPI_M_PC_INTERNAL_17 <= cpi_m_pc(18);
CPI_M_PC_INTERNAL_18 <= cpi_m_pc(19);
CPI_M_PC_INTERNAL_19 <= cpi_m_pc(20);
CPI_M_PC_INTERNAL_20 <= cpi_m_pc(21);
CPI_M_PC_INTERNAL_21 <= cpi_m_pc(22);
CPI_M_PC_INTERNAL_22 <= cpi_m_pc(23);
CPI_M_PC_INTERNAL_23 <= cpi_m_pc(24);
CPI_M_PC_INTERNAL_24 <= cpi_m_pc(25);
CPI_M_PC_INTERNAL_25 <= cpi_m_pc(26);
CPI_M_PC_INTERNAL_26 <= cpi_m_pc(27);
CPI_M_PC_INTERNAL_27 <= cpi_m_pc(28);
CPI_M_PC_INTERNAL_28 <= cpi_m_pc(29);
CPI_M_PC_INTERNAL_29 <= cpi_m_pc(30);
CPI_M_PC_INTERNAL_30 <= cpi_m_pc(31);
CPI_M_INST_INTERNAL <= cpi_m_inst(0);
CPI_M_INST_INTERNAL_0 <= cpi_m_inst(1);
CPI_M_INST_INTERNAL_1 <= cpi_m_inst(2);
CPI_M_INST_INTERNAL_2 <= cpi_m_inst(3);
CPI_M_INST_INTERNAL_3 <= cpi_m_inst(4);
CPI_M_INST_INTERNAL_4 <= cpi_m_inst(5);
CPI_M_INST_INTERNAL_5 <= cpi_m_inst(6);
CPI_M_INST_INTERNAL_6 <= cpi_m_inst(7);
CPI_M_INST_INTERNAL_7 <= cpi_m_inst(8);
CPI_M_INST_INTERNAL_8 <= cpi_m_inst(9);
CPI_M_INST_INTERNAL_9 <= cpi_m_inst(10);
CPI_M_INST_INTERNAL_10 <= cpi_m_inst(11);
CPI_M_INST_INTERNAL_11 <= cpi_m_inst(12);
CPI_M_INST_INTERNAL_12 <= cpi_m_inst(13);
CPI_M_INST_INTERNAL_13 <= cpi_m_inst(14);
CPI_M_INST_INTERNAL_14 <= cpi_m_inst(15);
CPI_M_INST_INTERNAL_15 <= cpi_m_inst(16);
CPI_M_INST_INTERNAL_16 <= cpi_m_inst(17);
CPI_M_INST_INTERNAL_17 <= cpi_m_inst(18);
CPI_M_INST_INTERNAL_18 <= cpi_m_inst(19);
CPI_M_INST_INTERNAL_19 <= cpi_m_inst(20);
CPI_M_INST_INTERNAL_20 <= cpi_m_inst(21);
CPI_M_INST_INTERNAL_21 <= cpi_m_inst(22);
CPI_M_INST_INTERNAL_22 <= cpi_m_inst(23);
CPI_M_INST_INTERNAL_23 <= cpi_m_inst(24);
CPI_M_INST_INTERNAL_24 <= cpi_m_inst(25);
CPI_M_INST_INTERNAL_25 <= cpi_m_inst(26);
CPI_M_INST_INTERNAL_26 <= cpi_m_inst(27);
CPI_M_INST_INTERNAL_27 <= cpi_m_inst(28);
CPI_M_INST_INTERNAL_28 <= cpi_m_inst(29);
CPI_M_INST_INTERNAL_29 <= cpi_m_inst(30);
CPI_M_INST_INTERNAL_30 <= cpi_m_inst(31);
CPI_M_CNT_INTERNAL <= cpi_m_cnt(0);
CPI_M_CNT_INTERNAL_0 <= cpi_m_cnt(1);
CPI_M_TRAP_INTERNAL <= cpi_m_trap;
CPI_M_ANNUL_INTERNAL <= cpi_m_annul;
CPI_M_PV_INTERNAL <= cpi_m_pv;
CPI_X_PC_INTERNAL <= cpi_x_pc(0);
CPI_X_PC_INTERNAL_0 <= cpi_x_pc(1);
CPI_X_PC_INTERNAL_1 <= cpi_x_pc(2);
CPI_X_PC_INTERNAL_2 <= cpi_x_pc(3);
CPI_X_PC_INTERNAL_3 <= cpi_x_pc(4);
CPI_X_PC_INTERNAL_4 <= cpi_x_pc(5);
CPI_X_PC_INTERNAL_5 <= cpi_x_pc(6);
CPI_X_PC_INTERNAL_6 <= cpi_x_pc(7);
CPI_X_PC_INTERNAL_7 <= cpi_x_pc(8);
CPI_X_PC_INTERNAL_8 <= cpi_x_pc(9);
CPI_X_PC_INTERNAL_9 <= cpi_x_pc(10);
CPI_X_PC_INTERNAL_10 <= cpi_x_pc(11);
CPI_X_PC_INTERNAL_11 <= cpi_x_pc(12);
CPI_X_PC_INTERNAL_12 <= cpi_x_pc(13);
CPI_X_PC_INTERNAL_13 <= cpi_x_pc(14);
CPI_X_PC_INTERNAL_14 <= cpi_x_pc(15);
CPI_X_PC_INTERNAL_15 <= cpi_x_pc(16);
CPI_X_PC_INTERNAL_16 <= cpi_x_pc(17);
CPI_X_PC_INTERNAL_17 <= cpi_x_pc(18);
CPI_X_PC_INTERNAL_18 <= cpi_x_pc(19);
CPI_X_PC_INTERNAL_19 <= cpi_x_pc(20);
CPI_X_PC_INTERNAL_20 <= cpi_x_pc(21);
CPI_X_PC_INTERNAL_21 <= cpi_x_pc(22);
CPI_X_PC_INTERNAL_22 <= cpi_x_pc(23);
CPI_X_PC_INTERNAL_23 <= cpi_x_pc(24);
CPI_X_PC_INTERNAL_24 <= cpi_x_pc(25);
CPI_X_PC_INTERNAL_25 <= cpi_x_pc(26);
CPI_X_PC_INTERNAL_26 <= cpi_x_pc(27);
CPI_X_PC_INTERNAL_27 <= cpi_x_pc(28);
CPI_X_PC_INTERNAL_28 <= cpi_x_pc(29);
CPI_X_PC_INTERNAL_29 <= cpi_x_pc(30);
CPI_X_PC_INTERNAL_30 <= cpi_x_pc(31);
CPI_X_INST_INTERNAL <= cpi_x_inst(0);
CPI_X_INST_INTERNAL_0 <= cpi_x_inst(1);
CPI_X_INST_INTERNAL_1 <= cpi_x_inst(2);
CPI_X_INST_INTERNAL_2 <= cpi_x_inst(3);
CPI_X_INST_INTERNAL_3 <= cpi_x_inst(4);
CPI_X_INST_INTERNAL_4 <= cpi_x_inst(5);
CPI_X_INST_INTERNAL_5 <= cpi_x_inst(6);
CPI_X_INST_INTERNAL_6 <= cpi_x_inst(7);
CPI_X_INST_INTERNAL_7 <= cpi_x_inst(8);
CPI_X_INST_INTERNAL_8 <= cpi_x_inst(9);
CPI_X_INST_INTERNAL_9 <= cpi_x_inst(10);
CPI_X_INST_INTERNAL_10 <= cpi_x_inst(11);
CPI_X_INST_INTERNAL_11 <= cpi_x_inst(12);
CPI_X_INST_INTERNAL_12 <= cpi_x_inst(13);
CPI_X_INST_INTERNAL_13 <= cpi_x_inst(14);
CPI_X_INST_INTERNAL_14 <= cpi_x_inst(15);
CPI_X_INST_INTERNAL_15 <= cpi_x_inst(16);
CPI_X_INST_INTERNAL_16 <= cpi_x_inst(17);
CPI_X_INST_INTERNAL_17 <= cpi_x_inst(18);
CPI_X_INST_INTERNAL_18 <= cpi_x_inst(19);
CPI_X_INST_INTERNAL_19 <= cpi_x_inst(20);
CPI_X_INST_INTERNAL_20 <= cpi_x_inst(21);
CPI_X_INST_INTERNAL_21 <= cpi_x_inst(22);
CPI_X_INST_INTERNAL_22 <= cpi_x_inst(23);
CPI_X_INST_INTERNAL_23 <= cpi_x_inst(24);
CPI_X_INST_INTERNAL_24 <= cpi_x_inst(25);
CPI_X_INST_INTERNAL_25 <= cpi_x_inst(26);
CPI_X_INST_INTERNAL_26 <= cpi_x_inst(27);
CPI_X_INST_INTERNAL_27 <= cpi_x_inst(28);
CPI_X_INST_INTERNAL_28 <= cpi_x_inst(29);
CPI_X_INST_INTERNAL_29 <= cpi_x_inst(30);
CPI_X_INST_INTERNAL_30 <= cpi_x_inst(31);
CPI_X_CNT_INTERNAL <= cpi_x_cnt(0);
CPI_X_CNT_INTERNAL_0 <= cpi_x_cnt(1);
CPI_X_TRAP_INTERNAL <= cpi_x_trap;
CPI_X_ANNUL_INTERNAL <= cpi_x_annul;
CPI_X_PV_INTERNAL <= cpi_x_pv;
CPI_LDDATA_INTERNAL <= cpi_lddata(0);
CPI_LDDATA_INTERNAL_0 <= cpi_lddata(1);
CPI_LDDATA_INTERNAL_1 <= cpi_lddata(2);
CPI_LDDATA_INTERNAL_2 <= cpi_lddata(3);
CPI_LDDATA_INTERNAL_3 <= cpi_lddata(4);
CPI_LDDATA_INTERNAL_4 <= cpi_lddata(5);
CPI_LDDATA_INTERNAL_5 <= cpi_lddata(6);
CPI_LDDATA_INTERNAL_6 <= cpi_lddata(7);
CPI_LDDATA_INTERNAL_7 <= cpi_lddata(8);
CPI_LDDATA_INTERNAL_8 <= cpi_lddata(9);
CPI_LDDATA_INTERNAL_9 <= cpi_lddata(10);
CPI_LDDATA_INTERNAL_10 <= cpi_lddata(11);
CPI_LDDATA_INTERNAL_11 <= cpi_lddata(12);
CPI_LDDATA_INTERNAL_12 <= cpi_lddata(13);
CPI_LDDATA_INTERNAL_13 <= cpi_lddata(14);
CPI_LDDATA_INTERNAL_14 <= cpi_lddata(15);
CPI_LDDATA_INTERNAL_15 <= cpi_lddata(16);
CPI_LDDATA_INTERNAL_16 <= cpi_lddata(17);
CPI_LDDATA_INTERNAL_17 <= cpi_lddata(18);
CPI_LDDATA_INTERNAL_18 <= cpi_lddata(19);
CPI_LDDATA_INTERNAL_19 <= cpi_lddata(20);
CPI_LDDATA_INTERNAL_20 <= cpi_lddata(21);
CPI_LDDATA_INTERNAL_21 <= cpi_lddata(22);
CPI_LDDATA_INTERNAL_22 <= cpi_lddata(23);
CPI_LDDATA_INTERNAL_23 <= cpi_lddata(24);
CPI_LDDATA_INTERNAL_24 <= cpi_lddata(25);
CPI_LDDATA_INTERNAL_25 <= cpi_lddata(26);
CPI_LDDATA_INTERNAL_26 <= cpi_lddata(27);
CPI_LDDATA_INTERNAL_27 <= cpi_lddata(28);
CPI_LDDATA_INTERNAL_28 <= cpi_lddata(29);
CPI_LDDATA_INTERNAL_29 <= cpi_lddata(30);
CPI_LDDATA_INTERNAL_30 <= cpi_lddata(31);
CPI_DBG_ENABLE_INTERNAL <= cpi_dbg_enable;
CPI_DBG_WRITE_INTERNAL <= cpi_dbg_write;
CPI_DBG_FSR_INTERNAL <= cpi_dbg_fsr;
CPI_DBG_ADDR_INTERNAL <= cpi_dbg_addr(0);
CPI_DBG_ADDR_INTERNAL_0 <= cpi_dbg_addr(1);
CPI_DBG_ADDR_INTERNAL_1 <= cpi_dbg_addr(2);
CPI_DBG_ADDR_INTERNAL_2 <= cpi_dbg_addr(3);
CPI_DBG_ADDR_INTERNAL_3 <= cpi_dbg_addr(4);
CPI_DBG_DATA_INTERNAL <= cpi_dbg_data(0);
CPI_DBG_DATA_INTERNAL_0 <= cpi_dbg_data(1);
CPI_DBG_DATA_INTERNAL_1 <= cpi_dbg_data(2);
CPI_DBG_DATA_INTERNAL_2 <= cpi_dbg_data(3);
CPI_DBG_DATA_INTERNAL_3 <= cpi_dbg_data(4);
CPI_DBG_DATA_INTERNAL_4 <= cpi_dbg_data(5);
CPI_DBG_DATA_INTERNAL_5 <= cpi_dbg_data(6);
CPI_DBG_DATA_INTERNAL_6 <= cpi_dbg_data(7);
CPI_DBG_DATA_INTERNAL_7 <= cpi_dbg_data(8);
CPI_DBG_DATA_INTERNAL_8 <= cpi_dbg_data(9);
CPI_DBG_DATA_INTERNAL_9 <= cpi_dbg_data(10);
CPI_DBG_DATA_INTERNAL_10 <= cpi_dbg_data(11);
CPI_DBG_DATA_INTERNAL_11 <= cpi_dbg_data(12);
CPI_DBG_DATA_INTERNAL_12 <= cpi_dbg_data(13);
CPI_DBG_DATA_INTERNAL_13 <= cpi_dbg_data(14);
CPI_DBG_DATA_INTERNAL_14 <= cpi_dbg_data(15);
CPI_DBG_DATA_INTERNAL_15 <= cpi_dbg_data(16);
CPI_DBG_DATA_INTERNAL_16 <= cpi_dbg_data(17);
CPI_DBG_DATA_INTERNAL_17 <= cpi_dbg_data(18);
CPI_DBG_DATA_INTERNAL_18 <= cpi_dbg_data(19);
CPI_DBG_DATA_INTERNAL_19 <= cpi_dbg_data(20);
CPI_DBG_DATA_INTERNAL_20 <= cpi_dbg_data(21);
CPI_DBG_DATA_INTERNAL_21 <= cpi_dbg_data(22);
CPI_DBG_DATA_INTERNAL_22 <= cpi_dbg_data(23);
CPI_DBG_DATA_INTERNAL_23 <= cpi_dbg_data(24);
CPI_DBG_DATA_INTERNAL_24 <= cpi_dbg_data(25);
CPI_DBG_DATA_INTERNAL_25 <= cpi_dbg_data(26);
CPI_DBG_DATA_INTERNAL_26 <= cpi_dbg_data(27);
CPI_DBG_DATA_INTERNAL_27 <= cpi_dbg_data(28);
CPI_DBG_DATA_INTERNAL_28 <= cpi_dbg_data(29);
CPI_DBG_DATA_INTERNAL_29 <= cpi_dbg_data(30);
CPI_DBG_DATA_INTERNAL_30 <= cpi_dbg_data(31);
RFO1_DATA1_INTERNAL <= rfo1_data1(0);
RFO1_DATA1_INTERNAL_0 <= rfo1_data1(1);
RFO1_DATA1_INTERNAL_1 <= rfo1_data1(2);
RFO1_DATA1_INTERNAL_2 <= rfo1_data1(3);
RFO1_DATA1_INTERNAL_3 <= rfo1_data1(4);
RFO1_DATA1_INTERNAL_4 <= rfo1_data1(5);
RFO1_DATA1_INTERNAL_5 <= rfo1_data1(6);
RFO1_DATA1_INTERNAL_6 <= rfo1_data1(7);
RFO1_DATA1_INTERNAL_7 <= rfo1_data1(8);
RFO1_DATA1_INTERNAL_8 <= rfo1_data1(9);
RFO1_DATA1_INTERNAL_9 <= rfo1_data1(10);
RFO1_DATA1_INTERNAL_10 <= rfo1_data1(11);
RFO1_DATA1_INTERNAL_11 <= rfo1_data1(12);
RFO1_DATA1_INTERNAL_12 <= rfo1_data1(13);
RFO1_DATA1_INTERNAL_13 <= rfo1_data1(14);
RFO1_DATA1_INTERNAL_14 <= rfo1_data1(15);
RFO1_DATA1_INTERNAL_15 <= rfo1_data1(16);
RFO1_DATA1_INTERNAL_16 <= rfo1_data1(17);
RFO1_DATA1_INTERNAL_17 <= rfo1_data1(18);
RFO1_DATA1_INTERNAL_18 <= rfo1_data1(19);
RFO1_DATA1_INTERNAL_19 <= rfo1_data1(20);
RFO1_DATA1_INTERNAL_20 <= rfo1_data1(21);
RFO1_DATA1_INTERNAL_21 <= rfo1_data1(22);
RFO1_DATA1_INTERNAL_22 <= rfo1_data1(23);
RFO1_DATA1_INTERNAL_23 <= rfo1_data1(24);
RFO1_DATA1_INTERNAL_24 <= rfo1_data1(25);
RFO1_DATA1_INTERNAL_25 <= rfo1_data1(26);
RFO1_DATA1_INTERNAL_26 <= rfo1_data1(27);
RFO1_DATA1_INTERNAL_27 <= rfo1_data1(28);
RFO1_DATA1_INTERNAL_28 <= rfo1_data1(29);
RFO1_DATA1_INTERNAL_29 <= rfo1_data1(30);
RFO1_DATA1_INTERNAL_30 <= rfo1_data1(31);
RFO1_DATA2_INTERNAL <= rfo1_data2(0);
RFO1_DATA2_INTERNAL_0 <= rfo1_data2(1);
RFO1_DATA2_INTERNAL_1 <= rfo1_data2(2);
RFO1_DATA2_INTERNAL_2 <= rfo1_data2(3);
RFO1_DATA2_INTERNAL_3 <= rfo1_data2(4);
RFO1_DATA2_INTERNAL_4 <= rfo1_data2(5);
RFO1_DATA2_INTERNAL_5 <= rfo1_data2(6);
RFO1_DATA2_INTERNAL_6 <= rfo1_data2(7);
RFO1_DATA2_INTERNAL_7 <= rfo1_data2(8);
RFO1_DATA2_INTERNAL_8 <= rfo1_data2(9);
RFO1_DATA2_INTERNAL_9 <= rfo1_data2(10);
RFO1_DATA2_INTERNAL_10 <= rfo1_data2(11);
RFO1_DATA2_INTERNAL_11 <= rfo1_data2(12);
RFO1_DATA2_INTERNAL_12 <= rfo1_data2(13);
RFO1_DATA2_INTERNAL_13 <= rfo1_data2(14);
RFO1_DATA2_INTERNAL_14 <= rfo1_data2(15);
RFO1_DATA2_INTERNAL_15 <= rfo1_data2(16);
RFO1_DATA2_INTERNAL_16 <= rfo1_data2(17);
RFO1_DATA2_INTERNAL_17 <= rfo1_data2(18);
RFO1_DATA2_INTERNAL_18 <= rfo1_data2(19);
RFO1_DATA2_INTERNAL_19 <= rfo1_data2(20);
RFO1_DATA2_INTERNAL_20 <= rfo1_data2(21);
RFO1_DATA2_INTERNAL_21 <= rfo1_data2(22);
RFO1_DATA2_INTERNAL_22 <= rfo1_data2(23);
RFO1_DATA2_INTERNAL_23 <= rfo1_data2(24);
RFO1_DATA2_INTERNAL_24 <= rfo1_data2(25);
RFO1_DATA2_INTERNAL_25 <= rfo1_data2(26);
RFO1_DATA2_INTERNAL_26 <= rfo1_data2(27);
RFO1_DATA2_INTERNAL_27 <= rfo1_data2(28);
RFO1_DATA2_INTERNAL_28 <= rfo1_data2(29);
RFO1_DATA2_INTERNAL_29 <= rfo1_data2(30);
RFO1_DATA2_INTERNAL_30 <= rfo1_data2(31);
RFO2_DATA1_INTERNAL <= rfo2_data1(0);
RFO2_DATA1_INTERNAL_0 <= rfo2_data1(1);
RFO2_DATA1_INTERNAL_1 <= rfo2_data1(2);
RFO2_DATA1_INTERNAL_2 <= rfo2_data1(3);
RFO2_DATA1_INTERNAL_3 <= rfo2_data1(4);
RFO2_DATA1_INTERNAL_4 <= rfo2_data1(5);
RFO2_DATA1_INTERNAL_5 <= rfo2_data1(6);
RFO2_DATA1_INTERNAL_6 <= rfo2_data1(7);
RFO2_DATA1_INTERNAL_7 <= rfo2_data1(8);
RFO2_DATA1_INTERNAL_8 <= rfo2_data1(9);
RFO2_DATA1_INTERNAL_9 <= rfo2_data1(10);
RFO2_DATA1_INTERNAL_10 <= rfo2_data1(11);
RFO2_DATA1_INTERNAL_11 <= rfo2_data1(12);
RFO2_DATA1_INTERNAL_12 <= rfo2_data1(13);
RFO2_DATA1_INTERNAL_13 <= rfo2_data1(14);
RFO2_DATA1_INTERNAL_14 <= rfo2_data1(15);
RFO2_DATA1_INTERNAL_15 <= rfo2_data1(16);
RFO2_DATA1_INTERNAL_16 <= rfo2_data1(17);
RFO2_DATA1_INTERNAL_17 <= rfo2_data1(18);
RFO2_DATA1_INTERNAL_18 <= rfo2_data1(19);
RFO2_DATA1_INTERNAL_19 <= rfo2_data1(20);
RFO2_DATA1_INTERNAL_20 <= rfo2_data1(21);
RFO2_DATA1_INTERNAL_21 <= rfo2_data1(22);
RFO2_DATA1_INTERNAL_22 <= rfo2_data1(23);
RFO2_DATA1_INTERNAL_23 <= rfo2_data1(24);
RFO2_DATA1_INTERNAL_24 <= rfo2_data1(25);
RFO2_DATA1_INTERNAL_25 <= rfo2_data1(26);
RFO2_DATA1_INTERNAL_26 <= rfo2_data1(27);
RFO2_DATA1_INTERNAL_27 <= rfo2_data1(28);
RFO2_DATA1_INTERNAL_28 <= rfo2_data1(29);
RFO2_DATA1_INTERNAL_29 <= rfo2_data1(30);
RFO2_DATA1_INTERNAL_30 <= rfo2_data1(31);
RFO2_DATA2_INTERNAL <= rfo2_data2(0);
RFO2_DATA2_INTERNAL_0 <= rfo2_data2(1);
RFO2_DATA2_INTERNAL_1 <= rfo2_data2(2);
RFO2_DATA2_INTERNAL_2 <= rfo2_data2(3);
RFO2_DATA2_INTERNAL_3 <= rfo2_data2(4);
RFO2_DATA2_INTERNAL_4 <= rfo2_data2(5);
RFO2_DATA2_INTERNAL_5 <= rfo2_data2(6);
RFO2_DATA2_INTERNAL_6 <= rfo2_data2(7);
RFO2_DATA2_INTERNAL_7 <= rfo2_data2(8);
RFO2_DATA2_INTERNAL_8 <= rfo2_data2(9);
RFO2_DATA2_INTERNAL_9 <= rfo2_data2(10);
RFO2_DATA2_INTERNAL_10 <= rfo2_data2(11);
RFO2_DATA2_INTERNAL_11 <= rfo2_data2(12);
RFO2_DATA2_INTERNAL_12 <= rfo2_data2(13);
RFO2_DATA2_INTERNAL_13 <= rfo2_data2(14);
RFO2_DATA2_INTERNAL_14 <= rfo2_data2(15);
RFO2_DATA2_INTERNAL_15 <= rfo2_data2(16);
RFO2_DATA2_INTERNAL_16 <= rfo2_data2(17);
RFO2_DATA2_INTERNAL_17 <= rfo2_data2(18);
RFO2_DATA2_INTERNAL_18 <= rfo2_data2(19);
RFO2_DATA2_INTERNAL_19 <= rfo2_data2(20);
RFO2_DATA2_INTERNAL_20 <= rfo2_data2(21);
RFO2_DATA2_INTERNAL_21 <= rfo2_data2(22);
RFO2_DATA2_INTERNAL_22 <= rfo2_data2(23);
RFO2_DATA2_INTERNAL_23 <= rfo2_data2(24);
RFO2_DATA2_INTERNAL_24 <= rfo2_data2(25);
RFO2_DATA2_INTERNAL_25 <= rfo2_data2(26);
RFO2_DATA2_INTERNAL_26 <= rfo2_data2(27);
RFO2_DATA2_INTERNAL_27 <= rfo2_data2(28);
RFO2_DATA2_INTERNAL_28 <= rfo2_data2(29);
RFO2_DATA2_INTERNAL_29 <= rfo2_data2(30);
RFO2_DATA2_INTERNAL_30 <= rfo2_data2(31);
end beh;

