------------------------------------------------------------------------------
--  This file is a part of the GRLIB VHDL IP LIBRARY
--  Copyright (C) 2011, Aeroflex Gaisler AB - all rights reserved.
--
-- ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN 
-- ACCORDANCE WITH THE GAISLER LICENSE AGREEMENT AND MUST BE APPROVED 
-- IN ADVANCE IN WRITING.
------------------------------------------------------------------------------
--
-- Written by Synplicity
-- Product Version "E-2010.09"
-- Program "Synplify Pro", Mapper "maprc, Build 140R"
-- Mon Jan 31 16:02:13 2011
--

--
-- Written by Synplify Pro version Build 140R
-- Mon Jan 31 16:02:13 2011
--

--
library ieee, cycloneiii;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
--library synplify;
--use synplify.components.all;
use cycloneiii.cycloneiii_components.all;
library altera;
use altera.altera_primitives_components.all;

entity grlfpw_0_cycloneiii is
port(
  rst :  in std_logic;
  clk :  in std_logic;
  holdn :  in std_logic;
  cpi_flush :  in std_logic;
  cpi_exack :  in std_logic;
  cpi_a_rs1 : in std_logic_vector(4 downto 0);
  cpi_d_pc : in std_logic_vector(31 downto 0);
  cpi_d_inst : in std_logic_vector(31 downto 0);
  cpi_d_cnt : in std_logic_vector(1 downto 0);
  cpi_d_trap :  in std_logic;
  cpi_d_annul :  in std_logic;
  cpi_d_pv :  in std_logic;
  cpi_a_pc : in std_logic_vector(31 downto 0);
  cpi_a_inst : in std_logic_vector(31 downto 0);
  cpi_a_cnt : in std_logic_vector(1 downto 0);
  cpi_a_trap :  in std_logic;
  cpi_a_annul :  in std_logic;
  cpi_a_pv :  in std_logic;
  cpi_e_pc : in std_logic_vector(31 downto 0);
  cpi_e_inst : in std_logic_vector(31 downto 0);
  cpi_e_cnt : in std_logic_vector(1 downto 0);
  cpi_e_trap :  in std_logic;
  cpi_e_annul :  in std_logic;
  cpi_e_pv :  in std_logic;
  cpi_m_pc : in std_logic_vector(31 downto 0);
  cpi_m_inst : in std_logic_vector(31 downto 0);
  cpi_m_cnt : in std_logic_vector(1 downto 0);
  cpi_m_trap :  in std_logic;
  cpi_m_annul :  in std_logic;
  cpi_m_pv :  in std_logic;
  cpi_x_pc : in std_logic_vector(31 downto 0);
  cpi_x_inst : in std_logic_vector(31 downto 0);
  cpi_x_cnt : in std_logic_vector(1 downto 0);
  cpi_x_trap :  in std_logic;
  cpi_x_annul :  in std_logic;
  cpi_x_pv :  in std_logic;
  cpi_lddata : in std_logic_vector(31 downto 0);
  cpi_dbg_enable :  in std_logic;
  cpi_dbg_write :  in std_logic;
  cpi_dbg_fsr :  in std_logic;
  cpi_dbg_addr : in std_logic_vector(4 downto 0);
  cpi_dbg_data : in std_logic_vector(31 downto 0);
  cpo_data : out std_logic_vector(31 downto 0);
  cpo_exc :  out std_logic;
  cpo_cc : out std_logic_vector(1 downto 0);
  cpo_ccv :  out std_logic;
  cpo_ldlock :  out std_logic;
  cpo_holdn :  out std_logic;
  cpo_dbg_data : out std_logic_vector(31 downto 0);
  rfi1_rd1addr : out std_logic_vector(3 downto 0);
  rfi1_rd2addr : out std_logic_vector(3 downto 0);
  rfi1_wraddr : out std_logic_vector(3 downto 0);
  rfi1_wrdata : out std_logic_vector(31 downto 0);
  rfi1_ren1 :  out std_logic;
  rfi1_ren2 :  out std_logic;
  rfi1_wren :  out std_logic;
  rfi2_rd1addr : out std_logic_vector(3 downto 0);
  rfi2_rd2addr : out std_logic_vector(3 downto 0);
  rfi2_wraddr : out std_logic_vector(3 downto 0);
  rfi2_wrdata : out std_logic_vector(31 downto 0);
  rfi2_ren1 :  out std_logic;
  rfi2_ren2 :  out std_logic;
  rfi2_wren :  out std_logic;
  rfo1_data1 : in std_logic_vector(31 downto 0);
  rfo1_data2 : in std_logic_vector(31 downto 0);
  rfo2_data1 : in std_logic_vector(31 downto 0);
  rfo2_data2 : in std_logic_vector(31 downto 0));
end grlfpw_0_cycloneiii;

architecture beh of grlfpw_0_cycloneiii is
  signal devclrn : std_logic := '1';
  signal devpor : std_logic := '1';
  signal devoe : std_logic := '0';
  signal \GRLFPC2_0.FPI.OP2_X\ : std_logic_vector(63 downto 32);
  signal \GRLFPC2_0.R.FSR.RD\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\ : std_logic_vector(16 downto 0);
  signal \GRLFPC2_0.R.STATE\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.R.I.INST\ : std_logic_vector(31 downto 0);
  signal \GRLFPC2_0.R.FSR.TEM\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.R.I.EXC\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.R.FSR.AEXC\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.R.A.RS1\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.R.A.RS2\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.R.FSR.CEXC\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.R.FSR.FTT\ : std_logic_vector(2 downto 0);
  signal \GRLFPC2_0.R.I.RES\ : std_logic_vector(63 downto 0);
  signal \GRLFPC2_0.COMB.V.I.RES_1\ : std_logic_vector(63 to 63);
  signal \GRLFPC2_0.R.A.RF1REN\ : std_logic_vector(2 downto 1);
  signal \GRLFPC2_0.R.A.RF2REN\ : std_logic_vector(2 downto 1);
  signal \GRLFPC2_0.R.MK.LDOP_RET_1\ : std_logic_vector(8 downto 0);
  signal \GRLFPC2_0.R.MK.LDOP_RET_4\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.R.A.MOV_RET\ : std_logic_vector(15 downto 0);
  signal \GRLFPC2_0.R.A.SEQERR_RET_4\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.R.A.ST_RET_2\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.R.A.AFQ_RET\ : std_logic_vector(9 downto 5);
  signal \GRLFPC2_0.COMB.V.I.RES_6_X\ : std_logic_vector(63 to 63);
  signal \GRLFPC2_0.R.I.CC\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.R.I.PC_RET\ : std_logic_vector(29 downto 0);
  signal \GRLFPC2_0.R.I.PC_RET_30\ : std_logic_vector(29 downto 0);
  signal \GRLFPC2_0.R.I.EXC_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.COMB.RS1_1\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\ : std_logic_vector(31 downto 0);
  signal \GRLFPC2_0.COMB.V.E.STDATA_1_1\ : std_logic_vector(31 downto 0);
  signal \GRLFPC2_0.COMB.RF1REN_1_0_0\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.COMB.RS2_1\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.COMB.V.FSR.CEXC_1_1_X\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.COMB.V.FSR.CEXC_1_2\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.COMB.V.FSR.TEM_1_0_X\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.COMB.V.FSR.RD_1_0_X\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\ : std_logic_vector(85 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\ : std_logic_vector(377 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.MIXOIN\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\ : std_logic_vector(57 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\ : std_logic_vector(57 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_V\ : std_logic_vector(2 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\ : std_logic_vector(12 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\ : std_logic_vector(57 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\ : std_logic_vector(12 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\ : std_logic_vector(12 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL\ : std_logic_vector(8 downto 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_DIVMULTV\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_14\ : std_logic_vector(172 downto 141);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_1.SUM_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_50_1.SUM_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_X\ : std_logic_vector(83 downto 81);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\ : std_logic_vector(80 downto 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW\ : std_logic_vector(10 downto 8);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\ : std_logic_vector(57 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\ : std_logic_vector(57 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\ : std_logic_vector(257 downto 141);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\ : std_logic_vector(257 downto 245);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\ : std_logic_vector(57 downto 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN8_TEMP_U\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_3\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_33\ : std_logic_vector(244 downto 237);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\ : std_logic_vector(257 downto 250);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF_0\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\ : std_logic_vector(112 downto 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\ : std_logic_vector(112 downto 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_13_2\ : std_logic_vector(33 to 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_1\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.COMB.V.STATE_1_IV\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_1\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O18_0\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O2\ : std_logic_vector(59 downto 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\ : std_logic_vector(59 downto 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_16_1\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_10\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_6\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_5\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_7\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A18\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_14\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_8\ : std_logic_vector(36 to 36);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_O13\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_1_1\ : std_logic_vector(51 downto 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\ : std_logic_vector(61 downto 22);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\ : std_logic_vector(58 downto 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_2_1\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_2\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_3_1\ : std_logic_vector(36 to 36);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_16_2\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\ : std_logic_vector(48 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_1_1\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_5\ : std_logic_vector(57 downto 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\ : std_logic_vector(61 downto 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_1_1\ : std_logic_vector(62 to 62);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_7_1\ : std_logic_vector(34 to 34);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_15_3\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_15_4\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_18\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\ : std_logic_vector(50 downto 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A22_1\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_7_1\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_8_1\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_9_1\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_10_1\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_13_1\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_14_1\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_16_4\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_2\ : std_logic_vector(57 downto 7);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_5\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2\ : std_logic_vector(42 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12\ : std_logic_vector(26 to 26);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_14\ : std_logic_vector(34 downto 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_12\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1_A2\ : std_logic_vector(39 to 39);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_9\ : std_logic_vector(51 downto 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_7\ : std_logic_vector(62 to 62);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_2_0_I_O2\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_1\ : std_logic_vector(26 downto 17);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_0\ : std_logic_vector(53 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_12_I_O2\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12\ : std_logic_vector(44 downto 17);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_1\ : std_logic_vector(61 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_37\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_4\ : std_logic_vector(50 downto 7);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_4_1\ : std_logic_vector(50 to 50);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_11\ : std_logic_vector(62 downto 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_0\ : std_logic_vector(42 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_17\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_11_0_A2\ : std_logic_vector(19 to 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A26_1\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_36\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0_1\ : std_logic_vector(41 to 41);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_10_1_0_A2\ : std_logic_vector(53 to 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1_A2_1\ : std_logic_vector(39 to 39);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1_A2_1_1\ : std_logic_vector(39 to 39);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_14_0_A2\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_23\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_2\ : std_logic_vector(57 downto 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_0\ : std_logic_vector(29 downto 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_4_1\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_12_1\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\ : std_logic_vector(59 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_5\ : std_logic_vector(32 to 32);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A19_1\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_2_0\ : std_logic_vector(35 downto 25);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_3_0_O2\ : std_logic_vector(17 to 17);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_2_0_O2\ : std_logic_vector(17 to 17);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_2_A2_1\ : std_logic_vector(17 to 17);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_1\ : std_logic_vector(49 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_1\ : std_logic_vector(49 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_2\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_2\ : std_logic_vector(49 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3\ : std_logic_vector(49 to 49);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_12_1\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_12_1\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_9_1\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29\ : std_logic_vector(19 to 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\ : std_logic_vector(58 downto 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_16_1\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_1\ : std_logic_vector(58 downto 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_3\ : std_logic_vector(58 downto 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_5\ : std_logic_vector(58 downto 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A15_1\ : std_logic_vector(18 to 18);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A25_1\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_0\ : std_logic_vector(49 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0_1\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_8_1\ : std_logic_vector(34 to 34);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_9_1\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_2\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_13_1\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_6\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_2\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_23\ : std_logic_vector(53 to 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_0\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_7_1\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_O27_2\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A2_9\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_1\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_1_1\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_5\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_5_1\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_0\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_10_1\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_0_2\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_4_1\ : std_logic_vector(49 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_5_1\ : std_logic_vector(36 to 36);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_3\ : std_logic_vector(59 downto 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_1\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_5\ : std_logic_vector(59 downto 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_5_1\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_6\ : std_logic_vector(59 downto 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_3\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_6_2\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_1\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_4\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_1\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_1\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A28_1\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_14_1\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4\ : std_logic_vector(51 downto 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_1\ : std_logic_vector(51 downto 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A3\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_7\ : std_logic_vector(51 downto 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_5_1\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_7_2\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_0\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_5\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_6_1\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_2\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O21\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_1\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_1_2\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_4_2\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O13_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_6\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_5_3\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_4\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_4_2\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_2\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_2_1\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_1_2\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O18_4\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_2\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_2_1\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_1\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O18_6\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_0\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_12\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_11_2\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_10\ : std_logic_vector(49 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_9\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_4\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_4\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_14_2\ : std_logic_vector(59 downto 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_M16\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0\ : std_logic_vector(49 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_2\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_M2\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A3_3_2\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_3\ : std_logic_vector(29 downto 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X3\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_2_4\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_1\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A7_1\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O7_1\ : std_logic_vector(29 downto 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_13_1\ : std_logic_vector(34 to 34);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_12_2\ : std_logic_vector(34 to 34);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_6_1\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_7_2\ : std_logic_vector(34 to 34);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_5\ : std_logic_vector(34 to 34);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_4\ : std_logic_vector(34 to 34);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_2\ : std_logic_vector(34 to 34);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_1\ : std_logic_vector(34 to 34);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_M17\ : std_logic_vector(34 to 34);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O17_1\ : std_logic_vector(34 to 34);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A17_1\ : std_logic_vector(34 to 34);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_18\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_16\ : std_logic_vector(51 downto 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_14\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_13\ : std_logic_vector(51 downto 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_10_2\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_6\ : std_logic_vector(51 downto 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_5\ : std_logic_vector(51 downto 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\ : std_logic_vector(55 downto 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_4\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_3\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_3\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A21\ : std_logic_vector(51 downto 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A21_2\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_14\ : std_logic_vector(36 to 36);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_12\ : std_logic_vector(36 downto 32);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A13_1\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_7\ : std_logic_vector(36 downto 32);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_3\ : std_logic_vector(36 downto 32);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_2\ : std_logic_vector(36 downto 32);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_2_1\ : std_logic_vector(36 to 36);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_1\ : std_logic_vector(36 downto 32);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_0\ : std_logic_vector(36 to 36);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_0_2\ : std_logic_vector(36 to 36);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20\ : std_logic_vector(36 to 36);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_1_0\ : std_logic_vector(36 to 36);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_23\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_22\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_19\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_18\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_16\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_14\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_13\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_I_X2\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_13_1\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_10\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_9\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_8\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_7\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_3\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_2\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_I_A26_1\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_22\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_22_1\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_19\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_18_3\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_17\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_16\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_15\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_12\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_11\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_10\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_9\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_8\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_6\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_4\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_M2\ : std_logic_vector(59 downto 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_3\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_2_2\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_1\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O28_5\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A28\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_M2_0\ : std_logic_vector(57 downto 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_16_2\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_15\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_10\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_8\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_M21\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_2\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_2_2\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O21_2\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O21_3\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A21_1\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_22\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_18\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_17\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_16\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_15_2\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_13\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_16_1\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_11\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_8\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_7\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_6\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_4\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_3\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_2\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_O30_7\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_21_2\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_15\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_14\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_13\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A13\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_13_1\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_1\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_11\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_6\ : std_logic_vector(50 downto 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A19_2\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_8\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_6\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_5\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_4\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_2\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_0_2\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A19\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_4\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_24\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_24_3\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_23\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_21\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_19\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_17_1\ : std_logic_vector(52 downto 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_16\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_13\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_13_1\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_11\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_9\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_8\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_5\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_4\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_2\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O27_10\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_0\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A27\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_19\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_17\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_16\ : std_logic_vector(59 downto 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_15\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_14_3\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O23\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_12\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11\ : std_logic_vector(59 downto 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_10\ : std_logic_vector(59 downto 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_9\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_8_1\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_1\ : std_logic_vector(59 downto 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_0\ : std_logic_vector(59 downto 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_6\ : std_logic_vector(59 downto 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_20_2\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_18_1\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_17_2\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_13\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_10_1\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_7\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_6\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_4\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_3\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_X2_2\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_1\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_M24\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_O24_3\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_5_1\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_16_2\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_13_2\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_1\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_10\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_9\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_8\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_6\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_3\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_2\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_2_2\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_5\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O25\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_20\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_19\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_16\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_11\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_9\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_6\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_4\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_2\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_1\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_0\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A25\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_20_2\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_18_3\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_16_1\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_16\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_14\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_12\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_11\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_M27\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_8_2\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_7\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_6\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_X2_0\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_M27_0\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_2\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_1\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_O27_4\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_11_2\ : std_logic_vector(18 to 18);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_6\ : std_logic_vector(18 to 18);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_5\ : std_logic_vector(18 to 18);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_2\ : std_logic_vector(18 to 18);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_2_3\ : std_logic_vector(18 to 18);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_1\ : std_logic_vector(18 to 18);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_1_2\ : std_logic_vector(18 to 18);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_0\ : std_logic_vector(18 to 18);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_0\ : std_logic_vector(53 to 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_38\ : std_logic_vector(53 to 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_37\ : std_logic_vector(53 to 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_36\ : std_logic_vector(53 to 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_34_2\ : std_logic_vector(53 to 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_30\ : std_logic_vector(53 to 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_29\ : std_logic_vector(53 to 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_28\ : std_logic_vector(53 to 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_26_2\ : std_logic_vector(53 to 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_22\ : std_logic_vector(53 to 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_M22\ : std_logic_vector(53 to 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_21\ : std_logic_vector(53 to 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_9\ : std_logic_vector(53 to 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_20\ : std_logic_vector(53 to 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_11\ : std_logic_vector(53 to 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_21\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_12\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_11\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_9\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_8\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_7\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_5\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_4\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_M26\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_3\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O26_5\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_1\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_0\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O26_8\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A26\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O26_9\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_24\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_O28_5\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_22\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_19\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_17\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_16\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_15\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_14\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_11\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_O28_1\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_9\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_O28_6\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_4\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_3\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_M2_0\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_0\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_A28\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_20\ : std_logic_vector(52 to 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_20_4\ : std_logic_vector(52 to 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_12_2\ : std_logic_vector(52 to 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_18\ : std_logic_vector(52 downto 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11_1\ : std_logic_vector(52 to 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_8\ : std_logic_vector(52 to 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7\ : std_logic_vector(52 to 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7_1\ : std_logic_vector(52 to 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_4\ : std_logic_vector(52 to 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_5\ : std_logic_vector(52 to 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_2\ : std_logic_vector(52 downto 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_M23\ : std_logic_vector(52 to 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_8\ : std_logic_vector(52 downto 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_25\ : std_logic_vector(58 to 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_24\ : std_logic_vector(58 downto 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_23\ : std_logic_vector(58 to 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_22_1\ : std_logic_vector(58 to 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_21\ : std_logic_vector(58 downto 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_18\ : std_logic_vector(58 to 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_15\ : std_logic_vector(58 to 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_11\ : std_logic_vector(58 to 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_10\ : std_logic_vector(58 to 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_8\ : std_logic_vector(58 downto 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_7\ : std_logic_vector(58 downto 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_6\ : std_logic_vector(58 to 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_4\ : std_logic_vector(58 downto 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_0\ : std_logic_vector(58 downto 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O29_6\ : std_logic_vector(58 to 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_25_1\ : std_logic_vector(19 to 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_16\ : std_logic_vector(19 to 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_10_1\ : std_logic_vector(19 to 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_9\ : std_logic_vector(19 to 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_2\ : std_logic_vector(19 to 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_M2\ : std_logic_vector(19 to 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_M29\ : std_logic_vector(19 to 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_13\ : std_logic_vector(33 to 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7_2\ : std_logic_vector(33 to 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_7\ : std_logic_vector(33 to 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23\ : std_logic_vector(33 to 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_13\ : std_logic_vector(49 to 49);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_19\ : std_logic_vector(49 to 49);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_11\ : std_logic_vector(49 to 49);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_7\ : std_logic_vector(49 to 49);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_6\ : std_logic_vector(49 to 49);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O16\ : std_logic_vector(49 to 49);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A16\ : std_logic_vector(49 to 49);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_1\ : std_logic_vector(49 to 49);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_6\ : std_logic_vector(62 to 62);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_1_0_A2\ : std_logic_vector(25 to 25);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_3_I_O2\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_0_A2\ : std_logic_vector(46 downto 41);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_A26_17_0_A2\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_0_A2\ : std_logic_vector(15 to 15);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_0_0_A2\ : std_logic_vector(17 to 17);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_7\ : std_logic_vector(62 downto 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2\ : std_logic_vector(43 downto 10);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1_A2_0\ : std_logic_vector(39 to 39);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1\ : std_logic_vector(22 downto 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_1\ : std_logic_vector(38 to 38);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_4_0_A2\ : std_logic_vector(17 to 17);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_2\ : std_logic_vector(44 downto 35);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0\ : std_logic_vector(26 downto 17);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_0_A2\ : std_logic_vector(44 downto 28);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_0_A2_0\ : std_logic_vector(44 downto 28);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_17_1_I_O2\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O6_3\ : std_logic_vector(30 to 30);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O6_2\ : std_logic_vector(30 to 30);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O6_1\ : std_logic_vector(30 to 30);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A6_2\ : std_logic_vector(30 to 30);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A6_3\ : std_logic_vector(30 to 30);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O6\ : std_logic_vector(30 to 30);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A20\ : std_logic_vector(32 to 32);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O20_6\ : std_logic_vector(32 to 32);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O20_5\ : std_logic_vector(32 to 32);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O20_3\ : std_logic_vector(32 to 32);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_4\ : std_logic_vector(32 to 32);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_6\ : std_logic_vector(32 to 32);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_13\ : std_logic_vector(32 to 32);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_17\ : std_logic_vector(32 to 32);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A7\ : std_logic_vector(29 to 29);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O7_2\ : std_logic_vector(29 to 29);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O7_0\ : std_logic_vector(29 to 29);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_4\ : std_logic_vector(29 to 29);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_5\ : std_logic_vector(25 to 25);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_5_1\ : std_logic_vector(25 to 25);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_27\ : std_logic_vector(57 downto 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_2\ : std_logic_vector(25 to 25);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_A28_11_0_A2\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_26\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_2\ : std_logic_vector(17 to 17);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_3\ : std_logic_vector(17 to 17);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_10\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_20\ : std_logic_vector(34 to 34);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_O2_2\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_1\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A2_7\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_O2_3\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_M2\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_35\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_0_0_O2\ : std_logic_vector(34 to 34);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_6_I_O2\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1_A2_3\ : std_logic_vector(39 to 39);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_25\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_45\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_11_0_A2\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_30\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_A2_1\ : std_logic_vector(26 to 26);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_22\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_8_0_A2\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_5_0_A2\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\ : std_logic_vector(56 downto 10);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\ : std_logic_vector(54 downto 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\ : std_logic_vector(57 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\ : std_logic_vector(57 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\ : std_logic_vector(57 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\ : std_logic_vector(57 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\ : std_logic_vector(22 downto 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\ : std_logic_vector(115 downto 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\ : std_logic_vector(115 downto 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\ : std_logic_vector(257 downto 232);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS\ : std_logic_vector(9 downto 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0\ : std_logic_vector(236 downto 232);
  signal \GRLFPC2_0.COMB.RS1_1_0_X\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.COMB.RF2REN_1_0\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.COMB.RS1_1_1_X\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2_1\ : std_logic_vector(9 to 9);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.EXPYBUS_0\ : std_logic_vector(9 downto 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_1\ : std_logic_vector(7 to 7);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_2\ : std_logic_vector(9 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M14\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M2\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M11\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M8\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\ : std_logic_vector(57 downto 0);
  signal \GRLFPC2_0.COMB.DBGDATA_4_0_X\ : std_logic_vector(31 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\ : std_logic_vector(57 downto 1);
  signal \GRLFPC2_0.FPI.OP1_X\ : std_logic_vector(63 downto 32);
  signal \GRLFPC2_0.COMB.V.STATE_7_IV_I\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.COMB.V.I.PC_1\ : std_logic_vector(31 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_U\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_0\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\ : std_logic_vector(57 downto 8);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\ : std_logic_vector(114 downto 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\ : std_logic_vector(55 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\ : std_logic_vector(55 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\ : std_logic_vector(57 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\ : std_logic_vector(55 downto 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\ : std_logic_vector(57 downto 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\ : std_logic_vector(8 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\ : std_logic_vector(56 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP_2\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\ : std_logic_vector(8 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_2\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_1\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.WQSCTRL_0\ : std_logic_vector(67 to 67);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN8_TEMP_2\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1\ : std_logic_vector(51 downto 30);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.WQSCTRL\ : std_logic_vector(68 to 68);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_I_M\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.EXCEP_1_TZ\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.COMB.V.A.RF2REN_1\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.COMB.V.A.RF1REN_1\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.COMB.RF1REN_1_0_X\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.COMB.V.FSR.FCC_1_0_X\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.COMB.V.FSR.FCC_1_1_X\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.COMB.V.FSR.AEXC_6_I_M\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.U_RDN_1\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.COMB.WRADDR_5_M\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\ : std_logic_vector(56 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_0\ : std_logic_vector(57 downto 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS_2\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1_X\ : std_logic_vector(25 downto 23);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_T_3\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.COMB.WRDATA_4_X\ : std_logic_vector(62 downto 0);
  signal \GRLFPC2_0.WRDATA_0_X\ : std_logic_vector(63 downto 0);
  signal \GRLFPC2_0.COMB.RF2REN_1_0_X\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.COMB.WRADDR_5_X\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.COMB.WRADDR_5_I_M2_X\ : std_logic_vector(3 downto 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58_0\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.SELECTQUOBITS.NOTDIVC\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLBREGXZ.XZBREGLC_2\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_0\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.EXPYBUS\ : std_logic_vector(6 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_7_0\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_17_1\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_7_1\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_1_TZ\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_22_0\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_1_0_0\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_9_TZ\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_YY\ : std_logic_vector(10 downto 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX\ : std_logic_vector(7 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_9_0\ : std_logic_vector(34 to 34);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_12_0\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_18_1_0\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_4_1\ : std_logic_vector(59 downto 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_11_0\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_1_1_0\ : std_logic_vector(62 to 62);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_9_0\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_14_0\ : std_logic_vector(52 to 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_8_1\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_5_1\ : std_logic_vector(62 to 62);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_0\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_15_1\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_9_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_6_0\ : std_logic_vector(19 to 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_6_1\ : std_logic_vector(49 to 49);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7_0\ : std_logic_vector(59 downto 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_17_0\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A13_0\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_0_0\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A15_0\ : std_logic_vector(18 to 18);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_1_0\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_IV\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_3_1_0\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_3_TZ\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_4\ : std_logic_vector(6 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_5\ : std_logic_vector(6 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13_0\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_6_0\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_3_0\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_6_0\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_O2_1_0\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_2_1\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_8_0\ : std_logic_vector(51 downto 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_10_0\ : std_logic_vector(34 to 34);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_19_0\ : std_logic_vector(58 to 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_20_1_0\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_12_0\ : std_logic_vector(51 downto 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_5_0\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_13_1\ : std_logic_vector(52 to 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_21_1\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_11_0\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_14_0\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_4_0\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_27_1\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_22_1\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_0_0\ : std_logic_vector(62 to 62);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_0_1\ : std_logic_vector(62 to 62);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_21_0\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_8_1\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_11_0\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_11_1_0\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_20_0\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_18_1\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_3_0\ : std_logic_vector(18 to 18);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_3_1\ : std_logic_vector(18 to 18);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_9_0\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_9_1\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_4_0\ : std_logic_vector(31 to 31);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_4_0\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_10_0\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_24_1\ : std_logic_vector(53 to 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_20_0\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_6_1\ : std_logic_vector(33 to 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_17_1_0\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_3_1_0\ : std_logic_vector(34 to 34);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_10_0\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_16_0\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_12_0_0\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_9_1\ : std_logic_vector(49 to 49);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_8_1\ : std_logic_vector(49 to 49);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_17_0\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_17_1\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_0\ : std_logic_vector(49 to 49);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_3_0\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_5_0\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_16_0\ : std_logic_vector(36 to 36);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_16_1\ : std_logic_vector(36 to 36);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_0_0\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_10_1\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_2_0\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_5_0\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_25_0\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_25_1\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O29_1_0\ : std_logic_vector(58 to 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_10_0\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_11_0\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_15_0\ : std_logic_vector(36 to 36);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_10_1\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_9_0\ : std_logic_vector(18 to 18);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_1_0\ : std_logic_vector(50 downto 10);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_2_0\ : std_logic_vector(36 to 36);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_7_1_0\ : std_logic_vector(27 to 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0_0\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_6_0\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0_2\ : std_logic_vector(50 to 50);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_4_0\ : std_logic_vector(25 to 25);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_15_0\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_2_1\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_10_1\ : std_logic_vector(32 to 32);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_11_0\ : std_logic_vector(18 to 18);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_16_1\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0_1_0\ : std_logic_vector(51 to 51);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_2_1\ : std_logic_vector(58 to 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_5_0\ : std_logic_vector(59 downto 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_6_1\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_0_1\ : std_logic_vector(26 to 26);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_12_0\ : std_logic_vector(19 to 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_3_1\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_23_0\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_5_0\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_11_0\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_23_0\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_1_0\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.COMB.RF1REN_1_0_0_A2_1\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A6_2_1\ : std_logic_vector(30 to 30);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11_0\ : std_logic_vector(33 to 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_3_1\ : std_logic_vector(54 to 54);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_2_2\ : std_logic_vector(62 to 62);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_2_3\ : std_logic_vector(62 to 62);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_2_0\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_5_0\ : std_logic_vector(19 to 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_1_1\ : std_logic_vector(19 to 19);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_7_0\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_5_2\ : std_logic_vector(57 to 57);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0_0\ : std_logic_vector(43 downto 10);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_16_1\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_13_0\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_0_0\ : std_logic_vector(18 to 18);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_9_0\ : std_logic_vector(33 to 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_3_1\ : std_logic_vector(58 to 58);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_6_0\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_10_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_5_0\ : std_logic_vector(36 to 36);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_7_0\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_0_1\ : std_logic_vector(33 to 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_1_1\ : std_logic_vector(49 to 49);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_0_1\ : std_logic_vector(29 downto 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_9_3\ : std_logic_vector(52 to 52);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_2_2\ : std_logic_vector(59 to 59);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_2_0\ : std_logic_vector(50 to 50);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A22_0\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.EXTEND.TEMP_1\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A7_0\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW_0\ : std_logic_vector(77 to 77);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_1_0\ : std_logic_vector(38 to 38);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_0\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_2_0_O2_0\ : std_logic_vector(17 to 17);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1\ : std_logic_vector(26 to 26);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_1\ : std_logic_vector(22 to 22);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_0\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_1\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_2\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_3_0\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_5\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_6\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_8\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_9\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_11\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_13\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_14\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_17\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_19\ : std_logic_vector(11 to 11);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_0\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_1\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_6\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_7\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_10\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_12\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_13\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_14\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_15\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_16\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_17\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_18\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_23\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_0\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_7\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_10\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_12\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_14\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_16\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_18\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_19\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_20\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_21\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV_0\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_IV_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_1_0\ : std_logic_vector(5 to 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_9_0_A2\ : std_logic_vector(61 to 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_O2\ : std_logic_vector(25 to 25);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11_2\ : std_logic_vector(33 to 33);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_4_2\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_12\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_26_2\ : std_logic_vector(60 to 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_18_2\ : std_logic_vector(48 to 48);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_14_2\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_1_0_A2\ : std_logic_vector(62 to 62);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_0_I_O2\ : std_logic_vector(53 to 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_2_0_A2\ : std_logic_vector(55 to 55);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_12_0_A2\ : std_logic_vector(62 to 62);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW\ : std_logic_vector(77 to 77);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\ : std_logic_vector(113 downto 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\ : std_logic_vector(44 downto 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\ : std_logic_vector(55 downto 17);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_0_A\ : std_logic_vector(57 downto 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3_A\ : std_logic_vector(3 downto 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_A\ : std_logic_vector(54 downto 9);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3_A\ : std_logic_vector(9 downto 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0_A\ : std_logic_vector(35 downto 22);
  signal \GRLFPC2_0.COMB.V.FSR.CEXC_1_2_A_X\ : std_logic_vector(4 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM_A\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_14_A\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8_A\ : std_logic_vector(42 downto 10);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_A\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_19_A\ : std_logic_vector(47 to 47);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_A\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_IV_0_A\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4_A\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_0_S\ : std_logic_vector(56 to 56);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP1\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP2\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\ : std_logic_vector(85 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\ : std_logic_vector(15 downto 10);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\ : std_logic_vector(19 downto 8);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\ : std_logic_vector(231 downto 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_X_RETO\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\ : std_logic_vector(84 downto 53);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_RETO\ : std_logic_vector(6 downto 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_M_RETO\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\ : std_logic_vector(3 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_U_RETO\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO\ : std_logic_vector(4 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO\ : std_logic_vector(2 to 2);
  signal CPI_D_INST_RETO : std_logic_vector(12 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO\ : std_logic_vector(79 to 79);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M\ : std_logic_vector(4 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP2_RETI\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.EXTEND.TEMP_1_A_RETI\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN8_TEMP_2_A_RETI\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.EXTEND.TEMP_1_RETI\ : std_logic_vector(1 to 1);
  signal RFO2_DATA1_RETO : std_logic_vector(28 downto 27);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\ : std_logic_vector(85 downto 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\ : std_logic_vector(113 downto 60);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\ : std_logic_vector(85 downto 84);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM_A_RETI\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M11_RETI\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M2_RETI\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M8_RETI\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5_RETI\ : std_logic_vector(1 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13_RETI\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12_RETI\ : std_logic_vector(3 downto 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13_0_RETI\ : std_logic_vector(3 to 3);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2_RETO\ : std_logic_vector(13 to 13);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_7_1_RETO\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_RETO\ : std_logic_vector(6 downto 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1I\ : std_logic_vector(16 to 16);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS_2_RETI\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_RETI\ : std_logic_vector(16 downto 8);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS_RETI\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0_RETI\ : std_logic_vector(8 downto 5);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN8_TEMP_2_RETI\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122_RETI\ : std_logic_vector(4 to 4);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M14_RETI\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\ : std_logic_vector(77 downto 61);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2_1_RETI\ : std_logic_vector(9 to 9);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\ : std_logic_vector(3 downto 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\ : std_logic_vector(3 downto 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\ : std_logic_vector(1 to 1);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP1\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP2\ : std_logic_vector(2 to 2);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP1\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP2\ : std_logic_vector(0 to 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\ : std_logic_vector(6 to 6);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\ : std_logic_vector(85 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP2\ : std_logic_vector(15 to 15);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\ : std_logic_vector(85 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\ : std_logic_vector(85 downto 0);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\ : std_logic_vector(85 downto 78);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\ : std_logic_vector(85 downto 78);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\ : std_logic_vector(85 downto 78);
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\ : std_logic_vector(85 downto 78);
  signal CPO_DATAZ : std_logic_vector(31 downto 0);
  signal CPO_CCZ : std_logic_vector(1 downto 0);
  signal CPO_DBG_DATAZ : std_logic_vector(31 downto 0);
  signal RFI1_WRDATAZ : std_logic_vector(31 downto 0);
  signal RFI2_RD1ADDRZ : std_logic_vector(3 downto 0);
  signal RFI2_RD2ADDRZ : std_logic_vector(3 downto 0);
  signal RFI2_WRADDRZ : std_logic_vector(3 downto 0);
  signal RFI2_WRDATAZ : std_logic_vector(31 downto 0);
  signal RST_INTERNAL : std_logic ;
  signal CLK_INTERNAL : std_logic ;
  signal CPI_FLUSH_INTERNAL : std_logic ;
  signal CPI_EXACK_INTERNAL : std_logic ;
  signal CPI_A_RS1_INTERNAL : std_logic ;
  signal CPI_A_RS1_INTERNAL_0 : std_logic ;
  signal CPI_A_RS1_INTERNAL_1 : std_logic ;
  signal CPI_A_RS1_INTERNAL_2 : std_logic ;
  signal CPI_A_RS1_INTERNAL_3 : std_logic ;
  signal CPI_D_PC_INTERNAL : std_logic ;
  signal CPI_D_PC_INTERNAL_0 : std_logic ;
  signal CPI_D_PC_INTERNAL_1 : std_logic ;
  signal CPI_D_PC_INTERNAL_2 : std_logic ;
  signal CPI_D_PC_INTERNAL_3 : std_logic ;
  signal CPI_D_PC_INTERNAL_4 : std_logic ;
  signal CPI_D_PC_INTERNAL_5 : std_logic ;
  signal CPI_D_PC_INTERNAL_6 : std_logic ;
  signal CPI_D_PC_INTERNAL_7 : std_logic ;
  signal CPI_D_PC_INTERNAL_8 : std_logic ;
  signal CPI_D_PC_INTERNAL_9 : std_logic ;
  signal CPI_D_PC_INTERNAL_10 : std_logic ;
  signal CPI_D_PC_INTERNAL_11 : std_logic ;
  signal CPI_D_PC_INTERNAL_12 : std_logic ;
  signal CPI_D_PC_INTERNAL_13 : std_logic ;
  signal CPI_D_PC_INTERNAL_14 : std_logic ;
  signal CPI_D_PC_INTERNAL_15 : std_logic ;
  signal CPI_D_PC_INTERNAL_16 : std_logic ;
  signal CPI_D_PC_INTERNAL_17 : std_logic ;
  signal CPI_D_PC_INTERNAL_18 : std_logic ;
  signal CPI_D_PC_INTERNAL_19 : std_logic ;
  signal CPI_D_PC_INTERNAL_20 : std_logic ;
  signal CPI_D_PC_INTERNAL_21 : std_logic ;
  signal CPI_D_PC_INTERNAL_22 : std_logic ;
  signal CPI_D_PC_INTERNAL_23 : std_logic ;
  signal CPI_D_PC_INTERNAL_24 : std_logic ;
  signal CPI_D_PC_INTERNAL_25 : std_logic ;
  signal CPI_D_PC_INTERNAL_26 : std_logic ;
  signal CPI_D_PC_INTERNAL_27 : std_logic ;
  signal CPI_D_PC_INTERNAL_28 : std_logic ;
  signal CPI_D_PC_INTERNAL_29 : std_logic ;
  signal CPI_D_PC_INTERNAL_30 : std_logic ;
  signal CPI_D_INST_INTERNAL : std_logic ;
  signal CPI_D_INST_INTERNAL_0 : std_logic ;
  signal CPI_D_INST_INTERNAL_1 : std_logic ;
  signal CPI_D_INST_INTERNAL_2 : std_logic ;
  signal CPI_D_INST_INTERNAL_3 : std_logic ;
  signal CPI_D_INST_INTERNAL_4 : std_logic ;
  signal CPI_D_INST_INTERNAL_5 : std_logic ;
  signal CPI_D_INST_INTERNAL_6 : std_logic ;
  signal CPI_D_INST_INTERNAL_7 : std_logic ;
  signal CPI_D_INST_INTERNAL_8 : std_logic ;
  signal CPI_D_INST_INTERNAL_9 : std_logic ;
  signal CPI_D_INST_INTERNAL_10 : std_logic ;
  signal CPI_D_INST_INTERNAL_11 : std_logic ;
  signal CPI_D_INST_INTERNAL_12 : std_logic ;
  signal CPI_D_INST_INTERNAL_13 : std_logic ;
  signal CPI_D_INST_INTERNAL_14 : std_logic ;
  signal CPI_D_INST_INTERNAL_15 : std_logic ;
  signal CPI_D_INST_INTERNAL_16 : std_logic ;
  signal CPI_D_INST_INTERNAL_17 : std_logic ;
  signal CPI_D_INST_INTERNAL_18 : std_logic ;
  signal CPI_D_INST_INTERNAL_19 : std_logic ;
  signal CPI_D_INST_INTERNAL_20 : std_logic ;
  signal CPI_D_INST_INTERNAL_21 : std_logic ;
  signal CPI_D_INST_INTERNAL_22 : std_logic ;
  signal CPI_D_INST_INTERNAL_23 : std_logic ;
  signal CPI_D_INST_INTERNAL_24 : std_logic ;
  signal CPI_D_INST_INTERNAL_25 : std_logic ;
  signal CPI_D_INST_INTERNAL_26 : std_logic ;
  signal CPI_D_INST_INTERNAL_27 : std_logic ;
  signal CPI_D_INST_INTERNAL_28 : std_logic ;
  signal CPI_D_INST_INTERNAL_29 : std_logic ;
  signal CPI_D_INST_INTERNAL_30 : std_logic ;
  signal CPI_D_CNT_INTERNAL : std_logic ;
  signal CPI_D_CNT_INTERNAL_0 : std_logic ;
  signal CPI_D_TRAP_INTERNAL : std_logic ;
  signal CPI_D_ANNUL_INTERNAL : std_logic ;
  signal CPI_D_PV_INTERNAL : std_logic ;
  signal CPI_A_PC_INTERNAL : std_logic ;
  signal CPI_A_PC_INTERNAL_0 : std_logic ;
  signal CPI_A_PC_INTERNAL_1 : std_logic ;
  signal CPI_A_PC_INTERNAL_2 : std_logic ;
  signal CPI_A_PC_INTERNAL_3 : std_logic ;
  signal CPI_A_PC_INTERNAL_4 : std_logic ;
  signal CPI_A_PC_INTERNAL_5 : std_logic ;
  signal CPI_A_PC_INTERNAL_6 : std_logic ;
  signal CPI_A_PC_INTERNAL_7 : std_logic ;
  signal CPI_A_PC_INTERNAL_8 : std_logic ;
  signal CPI_A_PC_INTERNAL_9 : std_logic ;
  signal CPI_A_PC_INTERNAL_10 : std_logic ;
  signal CPI_A_PC_INTERNAL_11 : std_logic ;
  signal CPI_A_PC_INTERNAL_12 : std_logic ;
  signal CPI_A_PC_INTERNAL_13 : std_logic ;
  signal CPI_A_PC_INTERNAL_14 : std_logic ;
  signal CPI_A_PC_INTERNAL_15 : std_logic ;
  signal CPI_A_PC_INTERNAL_16 : std_logic ;
  signal CPI_A_PC_INTERNAL_17 : std_logic ;
  signal CPI_A_PC_INTERNAL_18 : std_logic ;
  signal CPI_A_PC_INTERNAL_19 : std_logic ;
  signal CPI_A_PC_INTERNAL_20 : std_logic ;
  signal CPI_A_PC_INTERNAL_21 : std_logic ;
  signal CPI_A_PC_INTERNAL_22 : std_logic ;
  signal CPI_A_PC_INTERNAL_23 : std_logic ;
  signal CPI_A_PC_INTERNAL_24 : std_logic ;
  signal CPI_A_PC_INTERNAL_25 : std_logic ;
  signal CPI_A_PC_INTERNAL_26 : std_logic ;
  signal CPI_A_PC_INTERNAL_27 : std_logic ;
  signal CPI_A_PC_INTERNAL_28 : std_logic ;
  signal CPI_A_PC_INTERNAL_29 : std_logic ;
  signal CPI_A_PC_INTERNAL_30 : std_logic ;
  signal CPI_A_INST_INTERNAL : std_logic ;
  signal CPI_A_INST_INTERNAL_0 : std_logic ;
  signal CPI_A_INST_INTERNAL_1 : std_logic ;
  signal CPI_A_INST_INTERNAL_2 : std_logic ;
  signal CPI_A_INST_INTERNAL_3 : std_logic ;
  signal CPI_A_INST_INTERNAL_4 : std_logic ;
  signal CPI_A_INST_INTERNAL_5 : std_logic ;
  signal CPI_A_INST_INTERNAL_6 : std_logic ;
  signal CPI_A_INST_INTERNAL_7 : std_logic ;
  signal CPI_A_INST_INTERNAL_8 : std_logic ;
  signal CPI_A_INST_INTERNAL_9 : std_logic ;
  signal CPI_A_INST_INTERNAL_10 : std_logic ;
  signal CPI_A_INST_INTERNAL_11 : std_logic ;
  signal CPI_A_INST_INTERNAL_12 : std_logic ;
  signal CPI_A_INST_INTERNAL_13 : std_logic ;
  signal CPI_A_INST_INTERNAL_14 : std_logic ;
  signal CPI_A_INST_INTERNAL_15 : std_logic ;
  signal CPI_A_INST_INTERNAL_16 : std_logic ;
  signal CPI_A_INST_INTERNAL_17 : std_logic ;
  signal CPI_A_INST_INTERNAL_18 : std_logic ;
  signal CPI_A_INST_INTERNAL_19 : std_logic ;
  signal CPI_A_INST_INTERNAL_20 : std_logic ;
  signal CPI_A_INST_INTERNAL_21 : std_logic ;
  signal CPI_A_INST_INTERNAL_22 : std_logic ;
  signal CPI_A_INST_INTERNAL_23 : std_logic ;
  signal CPI_A_INST_INTERNAL_24 : std_logic ;
  signal CPI_A_INST_INTERNAL_25 : std_logic ;
  signal CPI_A_INST_INTERNAL_26 : std_logic ;
  signal CPI_A_INST_INTERNAL_27 : std_logic ;
  signal CPI_A_INST_INTERNAL_28 : std_logic ;
  signal CPI_A_INST_INTERNAL_29 : std_logic ;
  signal CPI_A_INST_INTERNAL_30 : std_logic ;
  signal CPI_A_CNT_INTERNAL : std_logic ;
  signal CPI_A_CNT_INTERNAL_0 : std_logic ;
  signal CPI_A_TRAP_INTERNAL : std_logic ;
  signal CPI_A_ANNUL_INTERNAL : std_logic ;
  signal CPI_A_PV_INTERNAL : std_logic ;
  signal CPI_E_PC_INTERNAL : std_logic ;
  signal CPI_E_PC_INTERNAL_0 : std_logic ;
  signal CPI_E_PC_INTERNAL_1 : std_logic ;
  signal CPI_E_PC_INTERNAL_2 : std_logic ;
  signal CPI_E_PC_INTERNAL_3 : std_logic ;
  signal CPI_E_PC_INTERNAL_4 : std_logic ;
  signal CPI_E_PC_INTERNAL_5 : std_logic ;
  signal CPI_E_PC_INTERNAL_6 : std_logic ;
  signal CPI_E_PC_INTERNAL_7 : std_logic ;
  signal CPI_E_PC_INTERNAL_8 : std_logic ;
  signal CPI_E_PC_INTERNAL_9 : std_logic ;
  signal CPI_E_PC_INTERNAL_10 : std_logic ;
  signal CPI_E_PC_INTERNAL_11 : std_logic ;
  signal CPI_E_PC_INTERNAL_12 : std_logic ;
  signal CPI_E_PC_INTERNAL_13 : std_logic ;
  signal CPI_E_PC_INTERNAL_14 : std_logic ;
  signal CPI_E_PC_INTERNAL_15 : std_logic ;
  signal CPI_E_PC_INTERNAL_16 : std_logic ;
  signal CPI_E_PC_INTERNAL_17 : std_logic ;
  signal CPI_E_PC_INTERNAL_18 : std_logic ;
  signal CPI_E_PC_INTERNAL_19 : std_logic ;
  signal CPI_E_PC_INTERNAL_20 : std_logic ;
  signal CPI_E_PC_INTERNAL_21 : std_logic ;
  signal CPI_E_PC_INTERNAL_22 : std_logic ;
  signal CPI_E_PC_INTERNAL_23 : std_logic ;
  signal CPI_E_PC_INTERNAL_24 : std_logic ;
  signal CPI_E_PC_INTERNAL_25 : std_logic ;
  signal CPI_E_PC_INTERNAL_26 : std_logic ;
  signal CPI_E_PC_INTERNAL_27 : std_logic ;
  signal CPI_E_PC_INTERNAL_28 : std_logic ;
  signal CPI_E_PC_INTERNAL_29 : std_logic ;
  signal CPI_E_PC_INTERNAL_30 : std_logic ;
  signal CPI_E_INST_INTERNAL : std_logic ;
  signal CPI_E_INST_INTERNAL_0 : std_logic ;
  signal CPI_E_INST_INTERNAL_1 : std_logic ;
  signal CPI_E_INST_INTERNAL_2 : std_logic ;
  signal CPI_E_INST_INTERNAL_3 : std_logic ;
  signal CPI_E_INST_INTERNAL_4 : std_logic ;
  signal CPI_E_INST_INTERNAL_5 : std_logic ;
  signal CPI_E_INST_INTERNAL_6 : std_logic ;
  signal CPI_E_INST_INTERNAL_7 : std_logic ;
  signal CPI_E_INST_INTERNAL_8 : std_logic ;
  signal CPI_E_INST_INTERNAL_9 : std_logic ;
  signal CPI_E_INST_INTERNAL_10 : std_logic ;
  signal CPI_E_INST_INTERNAL_11 : std_logic ;
  signal CPI_E_INST_INTERNAL_12 : std_logic ;
  signal CPI_E_INST_INTERNAL_13 : std_logic ;
  signal CPI_E_INST_INTERNAL_14 : std_logic ;
  signal CPI_E_INST_INTERNAL_15 : std_logic ;
  signal CPI_E_INST_INTERNAL_16 : std_logic ;
  signal CPI_E_INST_INTERNAL_17 : std_logic ;
  signal CPI_E_INST_INTERNAL_18 : std_logic ;
  signal CPI_E_INST_INTERNAL_19 : std_logic ;
  signal CPI_E_INST_INTERNAL_20 : std_logic ;
  signal CPI_E_INST_INTERNAL_21 : std_logic ;
  signal CPI_E_INST_INTERNAL_22 : std_logic ;
  signal CPI_E_INST_INTERNAL_23 : std_logic ;
  signal CPI_E_INST_INTERNAL_24 : std_logic ;
  signal CPI_E_INST_INTERNAL_25 : std_logic ;
  signal CPI_E_INST_INTERNAL_26 : std_logic ;
  signal CPI_E_INST_INTERNAL_27 : std_logic ;
  signal CPI_E_INST_INTERNAL_28 : std_logic ;
  signal CPI_E_INST_INTERNAL_29 : std_logic ;
  signal CPI_E_INST_INTERNAL_30 : std_logic ;
  signal CPI_E_CNT_INTERNAL : std_logic ;
  signal CPI_E_CNT_INTERNAL_0 : std_logic ;
  signal CPI_E_TRAP_INTERNAL : std_logic ;
  signal CPI_E_ANNUL_INTERNAL : std_logic ;
  signal CPI_E_PV_INTERNAL : std_logic ;
  signal CPI_M_PC_INTERNAL : std_logic ;
  signal CPI_M_PC_INTERNAL_0 : std_logic ;
  signal CPI_M_PC_INTERNAL_1 : std_logic ;
  signal CPI_M_PC_INTERNAL_2 : std_logic ;
  signal CPI_M_PC_INTERNAL_3 : std_logic ;
  signal CPI_M_PC_INTERNAL_4 : std_logic ;
  signal CPI_M_PC_INTERNAL_5 : std_logic ;
  signal CPI_M_PC_INTERNAL_6 : std_logic ;
  signal CPI_M_PC_INTERNAL_7 : std_logic ;
  signal CPI_M_PC_INTERNAL_8 : std_logic ;
  signal CPI_M_PC_INTERNAL_9 : std_logic ;
  signal CPI_M_PC_INTERNAL_10 : std_logic ;
  signal CPI_M_PC_INTERNAL_11 : std_logic ;
  signal CPI_M_PC_INTERNAL_12 : std_logic ;
  signal CPI_M_PC_INTERNAL_13 : std_logic ;
  signal CPI_M_PC_INTERNAL_14 : std_logic ;
  signal CPI_M_PC_INTERNAL_15 : std_logic ;
  signal CPI_M_PC_INTERNAL_16 : std_logic ;
  signal CPI_M_PC_INTERNAL_17 : std_logic ;
  signal CPI_M_PC_INTERNAL_18 : std_logic ;
  signal CPI_M_PC_INTERNAL_19 : std_logic ;
  signal CPI_M_PC_INTERNAL_20 : std_logic ;
  signal CPI_M_PC_INTERNAL_21 : std_logic ;
  signal CPI_M_PC_INTERNAL_22 : std_logic ;
  signal CPI_M_PC_INTERNAL_23 : std_logic ;
  signal CPI_M_PC_INTERNAL_24 : std_logic ;
  signal CPI_M_PC_INTERNAL_25 : std_logic ;
  signal CPI_M_PC_INTERNAL_26 : std_logic ;
  signal CPI_M_PC_INTERNAL_27 : std_logic ;
  signal CPI_M_PC_INTERNAL_28 : std_logic ;
  signal CPI_M_PC_INTERNAL_29 : std_logic ;
  signal CPI_M_PC_INTERNAL_30 : std_logic ;
  signal CPI_M_INST_INTERNAL : std_logic ;
  signal CPI_M_INST_INTERNAL_0 : std_logic ;
  signal CPI_M_INST_INTERNAL_1 : std_logic ;
  signal CPI_M_INST_INTERNAL_2 : std_logic ;
  signal CPI_M_INST_INTERNAL_3 : std_logic ;
  signal CPI_M_INST_INTERNAL_4 : std_logic ;
  signal CPI_M_INST_INTERNAL_5 : std_logic ;
  signal CPI_M_INST_INTERNAL_6 : std_logic ;
  signal CPI_M_INST_INTERNAL_7 : std_logic ;
  signal CPI_M_INST_INTERNAL_8 : std_logic ;
  signal CPI_M_INST_INTERNAL_9 : std_logic ;
  signal CPI_M_INST_INTERNAL_10 : std_logic ;
  signal CPI_M_INST_INTERNAL_11 : std_logic ;
  signal CPI_M_INST_INTERNAL_12 : std_logic ;
  signal CPI_M_INST_INTERNAL_13 : std_logic ;
  signal CPI_M_INST_INTERNAL_14 : std_logic ;
  signal CPI_M_INST_INTERNAL_15 : std_logic ;
  signal CPI_M_INST_INTERNAL_16 : std_logic ;
  signal CPI_M_INST_INTERNAL_17 : std_logic ;
  signal CPI_M_INST_INTERNAL_18 : std_logic ;
  signal CPI_M_INST_INTERNAL_19 : std_logic ;
  signal CPI_M_INST_INTERNAL_20 : std_logic ;
  signal CPI_M_INST_INTERNAL_21 : std_logic ;
  signal CPI_M_INST_INTERNAL_22 : std_logic ;
  signal CPI_M_INST_INTERNAL_23 : std_logic ;
  signal CPI_M_INST_INTERNAL_24 : std_logic ;
  signal CPI_M_INST_INTERNAL_25 : std_logic ;
  signal CPI_M_INST_INTERNAL_26 : std_logic ;
  signal CPI_M_INST_INTERNAL_27 : std_logic ;
  signal CPI_M_INST_INTERNAL_28 : std_logic ;
  signal CPI_M_INST_INTERNAL_29 : std_logic ;
  signal CPI_M_INST_INTERNAL_30 : std_logic ;
  signal CPI_M_CNT_INTERNAL : std_logic ;
  signal CPI_M_CNT_INTERNAL_0 : std_logic ;
  signal CPI_M_TRAP_INTERNAL : std_logic ;
  signal CPI_M_ANNUL_INTERNAL : std_logic ;
  signal CPI_M_PV_INTERNAL : std_logic ;
  signal CPI_X_PC_INTERNAL : std_logic ;
  signal CPI_X_PC_INTERNAL_0 : std_logic ;
  signal CPI_X_PC_INTERNAL_1 : std_logic ;
  signal CPI_X_PC_INTERNAL_2 : std_logic ;
  signal CPI_X_PC_INTERNAL_3 : std_logic ;
  signal CPI_X_PC_INTERNAL_4 : std_logic ;
  signal CPI_X_PC_INTERNAL_5 : std_logic ;
  signal CPI_X_PC_INTERNAL_6 : std_logic ;
  signal CPI_X_PC_INTERNAL_7 : std_logic ;
  signal CPI_X_PC_INTERNAL_8 : std_logic ;
  signal CPI_X_PC_INTERNAL_9 : std_logic ;
  signal CPI_X_PC_INTERNAL_10 : std_logic ;
  signal CPI_X_PC_INTERNAL_11 : std_logic ;
  signal CPI_X_PC_INTERNAL_12 : std_logic ;
  signal CPI_X_PC_INTERNAL_13 : std_logic ;
  signal CPI_X_PC_INTERNAL_14 : std_logic ;
  signal CPI_X_PC_INTERNAL_15 : std_logic ;
  signal CPI_X_PC_INTERNAL_16 : std_logic ;
  signal CPI_X_PC_INTERNAL_17 : std_logic ;
  signal CPI_X_PC_INTERNAL_18 : std_logic ;
  signal CPI_X_PC_INTERNAL_19 : std_logic ;
  signal CPI_X_PC_INTERNAL_20 : std_logic ;
  signal CPI_X_PC_INTERNAL_21 : std_logic ;
  signal CPI_X_PC_INTERNAL_22 : std_logic ;
  signal CPI_X_PC_INTERNAL_23 : std_logic ;
  signal CPI_X_PC_INTERNAL_24 : std_logic ;
  signal CPI_X_PC_INTERNAL_25 : std_logic ;
  signal CPI_X_PC_INTERNAL_26 : std_logic ;
  signal CPI_X_PC_INTERNAL_27 : std_logic ;
  signal CPI_X_PC_INTERNAL_28 : std_logic ;
  signal CPI_X_PC_INTERNAL_29 : std_logic ;
  signal CPI_X_PC_INTERNAL_30 : std_logic ;
  signal CPI_X_INST_INTERNAL : std_logic ;
  signal CPI_X_INST_INTERNAL_0 : std_logic ;
  signal CPI_X_INST_INTERNAL_1 : std_logic ;
  signal CPI_X_INST_INTERNAL_2 : std_logic ;
  signal CPI_X_INST_INTERNAL_3 : std_logic ;
  signal CPI_X_INST_INTERNAL_4 : std_logic ;
  signal CPI_X_INST_INTERNAL_5 : std_logic ;
  signal CPI_X_INST_INTERNAL_6 : std_logic ;
  signal CPI_X_INST_INTERNAL_7 : std_logic ;
  signal CPI_X_INST_INTERNAL_8 : std_logic ;
  signal CPI_X_INST_INTERNAL_9 : std_logic ;
  signal CPI_X_INST_INTERNAL_10 : std_logic ;
  signal CPI_X_INST_INTERNAL_11 : std_logic ;
  signal CPI_X_INST_INTERNAL_12 : std_logic ;
  signal CPI_X_INST_INTERNAL_13 : std_logic ;
  signal CPI_X_INST_INTERNAL_14 : std_logic ;
  signal CPI_X_INST_INTERNAL_15 : std_logic ;
  signal CPI_X_INST_INTERNAL_16 : std_logic ;
  signal CPI_X_INST_INTERNAL_17 : std_logic ;
  signal CPI_X_INST_INTERNAL_18 : std_logic ;
  signal CPI_X_INST_INTERNAL_19 : std_logic ;
  signal CPI_X_INST_INTERNAL_20 : std_logic ;
  signal CPI_X_INST_INTERNAL_21 : std_logic ;
  signal CPI_X_INST_INTERNAL_22 : std_logic ;
  signal CPI_X_INST_INTERNAL_23 : std_logic ;
  signal CPI_X_INST_INTERNAL_24 : std_logic ;
  signal CPI_X_INST_INTERNAL_25 : std_logic ;
  signal CPI_X_INST_INTERNAL_26 : std_logic ;
  signal CPI_X_INST_INTERNAL_27 : std_logic ;
  signal CPI_X_INST_INTERNAL_28 : std_logic ;
  signal CPI_X_INST_INTERNAL_29 : std_logic ;
  signal CPI_X_INST_INTERNAL_30 : std_logic ;
  signal CPI_X_CNT_INTERNAL : std_logic ;
  signal CPI_X_CNT_INTERNAL_0 : std_logic ;
  signal CPI_X_TRAP_INTERNAL : std_logic ;
  signal CPI_X_ANNUL_INTERNAL : std_logic ;
  signal CPI_X_PV_INTERNAL : std_logic ;
  signal CPI_LDDATA_INTERNAL : std_logic ;
  signal CPI_LDDATA_INTERNAL_0 : std_logic ;
  signal CPI_LDDATA_INTERNAL_1 : std_logic ;
  signal CPI_LDDATA_INTERNAL_2 : std_logic ;
  signal CPI_LDDATA_INTERNAL_3 : std_logic ;
  signal CPI_LDDATA_INTERNAL_4 : std_logic ;
  signal CPI_LDDATA_INTERNAL_5 : std_logic ;
  signal CPI_LDDATA_INTERNAL_6 : std_logic ;
  signal CPI_LDDATA_INTERNAL_7 : std_logic ;
  signal CPI_LDDATA_INTERNAL_8 : std_logic ;
  signal CPI_LDDATA_INTERNAL_9 : std_logic ;
  signal CPI_LDDATA_INTERNAL_10 : std_logic ;
  signal CPI_LDDATA_INTERNAL_11 : std_logic ;
  signal CPI_LDDATA_INTERNAL_12 : std_logic ;
  signal CPI_LDDATA_INTERNAL_13 : std_logic ;
  signal CPI_LDDATA_INTERNAL_14 : std_logic ;
  signal CPI_LDDATA_INTERNAL_15 : std_logic ;
  signal CPI_LDDATA_INTERNAL_16 : std_logic ;
  signal CPI_LDDATA_INTERNAL_17 : std_logic ;
  signal CPI_LDDATA_INTERNAL_18 : std_logic ;
  signal CPI_LDDATA_INTERNAL_19 : std_logic ;
  signal CPI_LDDATA_INTERNAL_20 : std_logic ;
  signal CPI_LDDATA_INTERNAL_21 : std_logic ;
  signal CPI_LDDATA_INTERNAL_22 : std_logic ;
  signal CPI_LDDATA_INTERNAL_23 : std_logic ;
  signal CPI_LDDATA_INTERNAL_24 : std_logic ;
  signal CPI_LDDATA_INTERNAL_25 : std_logic ;
  signal CPI_LDDATA_INTERNAL_26 : std_logic ;
  signal CPI_LDDATA_INTERNAL_27 : std_logic ;
  signal CPI_LDDATA_INTERNAL_28 : std_logic ;
  signal CPI_LDDATA_INTERNAL_29 : std_logic ;
  signal CPI_LDDATA_INTERNAL_30 : std_logic ;
  signal CPI_DBG_WRITE_INTERNAL : std_logic ;
  signal CPI_DBG_ADDR_INTERNAL_0 : std_logic ;
  signal CPI_DBG_ADDR_INTERNAL_1 : std_logic ;
  signal CPI_DBG_ADDR_INTERNAL_2 : std_logic ;
  signal CPI_DBG_ADDR_INTERNAL_3 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_0 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_1 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_2 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_3 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_4 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_5 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_6 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_7 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_8 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_9 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_10 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_11 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_12 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_13 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_14 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_15 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_16 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_17 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_18 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_19 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_20 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_21 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_22 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_23 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_24 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_25 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_26 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_27 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_28 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_29 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_30 : std_logic ;
  signal RFO1_DATA1_INTERNAL : std_logic ;
  signal RFO1_DATA1_INTERNAL_0 : std_logic ;
  signal RFO1_DATA1_INTERNAL_1 : std_logic ;
  signal RFO1_DATA1_INTERNAL_2 : std_logic ;
  signal RFO1_DATA1_INTERNAL_3 : std_logic ;
  signal RFO1_DATA1_INTERNAL_4 : std_logic ;
  signal RFO1_DATA1_INTERNAL_5 : std_logic ;
  signal RFO1_DATA1_INTERNAL_6 : std_logic ;
  signal RFO1_DATA1_INTERNAL_7 : std_logic ;
  signal RFO1_DATA1_INTERNAL_8 : std_logic ;
  signal RFO1_DATA1_INTERNAL_9 : std_logic ;
  signal RFO1_DATA1_INTERNAL_10 : std_logic ;
  signal RFO1_DATA1_INTERNAL_11 : std_logic ;
  signal RFO1_DATA1_INTERNAL_12 : std_logic ;
  signal RFO1_DATA1_INTERNAL_13 : std_logic ;
  signal RFO1_DATA1_INTERNAL_14 : std_logic ;
  signal RFO1_DATA1_INTERNAL_15 : std_logic ;
  signal RFO1_DATA1_INTERNAL_16 : std_logic ;
  signal RFO1_DATA1_INTERNAL_17 : std_logic ;
  signal RFO1_DATA1_INTERNAL_18 : std_logic ;
  signal RFO1_DATA1_INTERNAL_19 : std_logic ;
  signal RFO1_DATA1_INTERNAL_20 : std_logic ;
  signal RFO1_DATA1_INTERNAL_21 : std_logic ;
  signal RFO1_DATA1_INTERNAL_22 : std_logic ;
  signal RFO1_DATA1_INTERNAL_23 : std_logic ;
  signal RFO1_DATA1_INTERNAL_24 : std_logic ;
  signal RFO1_DATA1_INTERNAL_25 : std_logic ;
  signal RFO1_DATA1_INTERNAL_26 : std_logic ;
  signal RFO1_DATA1_INTERNAL_27 : std_logic ;
  signal RFO1_DATA1_INTERNAL_28 : std_logic ;
  signal RFO1_DATA1_INTERNAL_29 : std_logic ;
  signal RFO1_DATA1_INTERNAL_30 : std_logic ;
  signal RFO1_DATA2_INTERNAL : std_logic ;
  signal RFO1_DATA2_INTERNAL_0 : std_logic ;
  signal RFO1_DATA2_INTERNAL_1 : std_logic ;
  signal RFO1_DATA2_INTERNAL_2 : std_logic ;
  signal RFO1_DATA2_INTERNAL_3 : std_logic ;
  signal RFO1_DATA2_INTERNAL_4 : std_logic ;
  signal RFO1_DATA2_INTERNAL_5 : std_logic ;
  signal RFO1_DATA2_INTERNAL_6 : std_logic ;
  signal RFO1_DATA2_INTERNAL_7 : std_logic ;
  signal RFO1_DATA2_INTERNAL_8 : std_logic ;
  signal RFO1_DATA2_INTERNAL_9 : std_logic ;
  signal RFO1_DATA2_INTERNAL_10 : std_logic ;
  signal RFO1_DATA2_INTERNAL_11 : std_logic ;
  signal RFO1_DATA2_INTERNAL_12 : std_logic ;
  signal RFO1_DATA2_INTERNAL_13 : std_logic ;
  signal RFO1_DATA2_INTERNAL_14 : std_logic ;
  signal RFO1_DATA2_INTERNAL_15 : std_logic ;
  signal RFO1_DATA2_INTERNAL_16 : std_logic ;
  signal RFO1_DATA2_INTERNAL_17 : std_logic ;
  signal RFO1_DATA2_INTERNAL_18 : std_logic ;
  signal RFO1_DATA2_INTERNAL_19 : std_logic ;
  signal RFO1_DATA2_INTERNAL_20 : std_logic ;
  signal RFO1_DATA2_INTERNAL_21 : std_logic ;
  signal RFO1_DATA2_INTERNAL_22 : std_logic ;
  signal RFO1_DATA2_INTERNAL_23 : std_logic ;
  signal RFO1_DATA2_INTERNAL_24 : std_logic ;
  signal RFO1_DATA2_INTERNAL_25 : std_logic ;
  signal RFO1_DATA2_INTERNAL_26 : std_logic ;
  signal RFO1_DATA2_INTERNAL_27 : std_logic ;
  signal RFO1_DATA2_INTERNAL_28 : std_logic ;
  signal RFO1_DATA2_INTERNAL_29 : std_logic ;
  signal RFO1_DATA2_INTERNAL_30 : std_logic ;
  signal RFO2_DATA1_INTERNAL : std_logic ;
  signal RFO2_DATA1_INTERNAL_0 : std_logic ;
  signal RFO2_DATA1_INTERNAL_1 : std_logic ;
  signal RFO2_DATA1_INTERNAL_2 : std_logic ;
  signal RFO2_DATA1_INTERNAL_3 : std_logic ;
  signal RFO2_DATA1_INTERNAL_4 : std_logic ;
  signal RFO2_DATA1_INTERNAL_5 : std_logic ;
  signal RFO2_DATA1_INTERNAL_6 : std_logic ;
  signal RFO2_DATA1_INTERNAL_7 : std_logic ;
  signal RFO2_DATA1_INTERNAL_8 : std_logic ;
  signal RFO2_DATA1_INTERNAL_9 : std_logic ;
  signal RFO2_DATA1_INTERNAL_10 : std_logic ;
  signal RFO2_DATA1_INTERNAL_11 : std_logic ;
  signal RFO2_DATA1_INTERNAL_12 : std_logic ;
  signal RFO2_DATA1_INTERNAL_13 : std_logic ;
  signal RFO2_DATA1_INTERNAL_14 : std_logic ;
  signal RFO2_DATA1_INTERNAL_15 : std_logic ;
  signal RFO2_DATA1_INTERNAL_16 : std_logic ;
  signal RFO2_DATA1_INTERNAL_17 : std_logic ;
  signal RFO2_DATA1_INTERNAL_18 : std_logic ;
  signal RFO2_DATA1_INTERNAL_19 : std_logic ;
  signal RFO2_DATA1_INTERNAL_20 : std_logic ;
  signal RFO2_DATA1_INTERNAL_21 : std_logic ;
  signal RFO2_DATA1_INTERNAL_22 : std_logic ;
  signal RFO2_DATA1_INTERNAL_23 : std_logic ;
  signal RFO2_DATA1_INTERNAL_24 : std_logic ;
  signal RFO2_DATA1_INTERNAL_25 : std_logic ;
  signal RFO2_DATA1_INTERNAL_26 : std_logic ;
  signal RFO2_DATA1_INTERNAL_27 : std_logic ;
  signal RFO2_DATA1_INTERNAL_28 : std_logic ;
  signal RFO2_DATA1_INTERNAL_29 : std_logic ;
  signal RFO2_DATA1_INTERNAL_30 : std_logic ;
  signal RFO2_DATA2_INTERNAL : std_logic ;
  signal RFO2_DATA2_INTERNAL_0 : std_logic ;
  signal RFO2_DATA2_INTERNAL_1 : std_logic ;
  signal RFO2_DATA2_INTERNAL_2 : std_logic ;
  signal RFO2_DATA2_INTERNAL_3 : std_logic ;
  signal RFO2_DATA2_INTERNAL_4 : std_logic ;
  signal RFO2_DATA2_INTERNAL_5 : std_logic ;
  signal RFO2_DATA2_INTERNAL_6 : std_logic ;
  signal RFO2_DATA2_INTERNAL_7 : std_logic ;
  signal RFO2_DATA2_INTERNAL_8 : std_logic ;
  signal RFO2_DATA2_INTERNAL_9 : std_logic ;
  signal RFO2_DATA2_INTERNAL_10 : std_logic ;
  signal RFO2_DATA2_INTERNAL_11 : std_logic ;
  signal RFO2_DATA2_INTERNAL_12 : std_logic ;
  signal RFO2_DATA2_INTERNAL_13 : std_logic ;
  signal RFO2_DATA2_INTERNAL_14 : std_logic ;
  signal RFO2_DATA2_INTERNAL_15 : std_logic ;
  signal RFO2_DATA2_INTERNAL_16 : std_logic ;
  signal RFO2_DATA2_INTERNAL_17 : std_logic ;
  signal RFO2_DATA2_INTERNAL_18 : std_logic ;
  signal RFO2_DATA2_INTERNAL_19 : std_logic ;
  signal RFO2_DATA2_INTERNAL_20 : std_logic ;
  signal RFO2_DATA2_INTERNAL_21 : std_logic ;
  signal RFO2_DATA2_INTERNAL_22 : std_logic ;
  signal RFO2_DATA2_INTERNAL_23 : std_logic ;
  signal RFO2_DATA2_INTERNAL_24 : std_logic ;
  signal RFO2_DATA2_INTERNAL_25 : std_logic ;
  signal RFO2_DATA2_INTERNAL_26 : std_logic ;
  signal RFO2_DATA2_INTERNAL_27 : std_logic ;
  signal RFO2_DATA2_INTERNAL_28 : std_logic ;
  signal RFO2_DATA2_INTERNAL_29 : std_logic ;
  signal RFO2_DATA2_INTERNAL_30 : std_logic ;
  signal VCC : std_logic ;
  signal GND : std_logic ;
  signal \GRLFPC2_0.FPI.START\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD16\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD18\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD19\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD20\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD21\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD22\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD23\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD24\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD25\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD26\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD27\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD28\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD29\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD30\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD31\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD32\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD33\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD34\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD35\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD36\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD37\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD38\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD39\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD40\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD41\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD42\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD43\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD44\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD45\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD46\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD47\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD48\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD49\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD50\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD51\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD52\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD53\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD54\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.SIGNRESULT\ : std_logic ;
  signal \GRLFPC2_0.R.I.EXEC\ : std_logic ;
  signal \GRLFPC2_0.R.X.LD\ : std_logic ;
  signal \GRLFPC2_0.R.X.AFSR\ : std_logic ;
  signal \GRLFPC2_0.R.X.SEQERR\ : std_logic ;
  signal \GRLFPC2_0.R.X.FPOP\ : std_logic ;
  signal \GRLFPC2_0.R.E.FPOP\ : std_logic ;
  signal \GRLFPC2_0.R.M.FPOP\ : std_logic ;
  signal \GRLFPC2_0.R.MK.HOLDN2\ : std_logic ;
  signal \GRLFPC2_0.R.I.V\ : std_logic ;
  signal \GRLFPC2_0.R.M.LD\ : std_logic ;
  signal \GRLFPC2_0.R.E.LD\ : std_logic ;
  signal \GRLFPC2_0.R.A.LD\ : std_logic ;
  signal \GRLFPC2_0.R.A.FPOP\ : std_logic ;
  signal \GRLFPC2_0.R.X.AFQ\ : std_logic ;
  signal \GRLFPC2_0.R.I.RDD\ : std_logic ;
  signal \GRLFPC2_0.R.X.RDD\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.NONSTD\ : std_logic ;
  signal \GRLFPC2_0.R.M.SEQERR\ : std_logic ;
  signal \GRLFPC2_0.R.A.RDD\ : std_logic ;
  signal \GRLFPC2_0.R.E.RDD\ : std_logic ;
  signal \GRLFPC2_0.R.M.RDD\ : std_logic ;
  signal \GRLFPC2_0.N_95\ : std_logic ;
  signal \GRLFPC2_0.N_96\ : std_logic ;
  signal \GRLFPC2_0.N_97\ : std_logic ;
  signal \GRLFPC2_0.N_98\ : std_logic ;
  signal \GRLFPC2_0.N_99\ : std_logic ;
  signal \GRLFPC2_0.N_100\ : std_logic ;
  signal \GRLFPC2_0.N_101\ : std_logic ;
  signal \GRLFPC2_0.N_102\ : std_logic ;
  signal \GRLFPC2_0.N_103\ : std_logic ;
  signal \GRLFPC2_0.N_104\ : std_logic ;
  signal \GRLFPC2_0.N_105\ : std_logic ;
  signal \GRLFPC2_0.N_106\ : std_logic ;
  signal \GRLFPC2_0.N_107\ : std_logic ;
  signal \GRLFPC2_0.N_108\ : std_logic ;
  signal \GRLFPC2_0.N_109\ : std_logic ;
  signal \GRLFPC2_0.N_110\ : std_logic ;
  signal \GRLFPC2_0.N_111\ : std_logic ;
  signal \GRLFPC2_0.N_112\ : std_logic ;
  signal \GRLFPC2_0.N_113\ : std_logic ;
  signal \GRLFPC2_0.N_114\ : std_logic ;
  signal \GRLFPC2_0.N_115\ : std_logic ;
  signal \GRLFPC2_0.N_116\ : std_logic ;
  signal \GRLFPC2_0.N_117\ : std_logic ;
  signal \GRLFPC2_0.N_118\ : std_logic ;
  signal \GRLFPC2_0.N_119\ : std_logic ;
  signal \GRLFPC2_0.N_120\ : std_logic ;
  signal \GRLFPC2_0.N_121\ : std_logic ;
  signal \GRLFPC2_0.N_122\ : std_logic ;
  signal \GRLFPC2_0.N_123\ : std_logic ;
  signal \GRLFPC2_0.N_124\ : std_logic ;
  signal \GRLFPC2_0.N_125\ : std_logic ;
  signal \GRLFPC2_0.N_126\ : std_logic ;
  signal \GRLFPC2_0.N_127\ : std_logic ;
  signal \GRLFPC2_0.N_128\ : std_logic ;
  signal \GRLFPC2_0.N_129\ : std_logic ;
  signal \GRLFPC2_0.N_130\ : std_logic ;
  signal \GRLFPC2_0.N_131\ : std_logic ;
  signal \GRLFPC2_0.N_132\ : std_logic ;
  signal \GRLFPC2_0.N_133\ : std_logic ;
  signal \GRLFPC2_0.N_134\ : std_logic ;
  signal \GRLFPC2_0.N_135\ : std_logic ;
  signal \GRLFPC2_0.N_136\ : std_logic ;
  signal \GRLFPC2_0.N_137\ : std_logic ;
  signal \GRLFPC2_0.R.MK.LDOP_RET\ : std_logic ;
  signal \GRLFPC2_0.R.MK.LDOP_RET_3\ : std_logic ;
  signal \GRLFPC2_0.R.MK.LDOP_RET_6\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.MK.RST_1_0_A2\ : std_logic ;
  signal \GRLFPC2_0.R.MK.RST2\ : std_logic ;
  signal \GRLFPC2_0.R.MK.RST_RET\ : std_logic ;
  signal \GRLFPC2_0.R.MK.RST_RET_6\ : std_logic ;
  signal \GRLFPC2_0.R.MK.BUSY_RET_4\ : std_logic ;
  signal \GRLFPC2_0.R.MK.RST_RET_2\ : std_logic ;
  signal \GRLFPC2_0.R.MK.BUSY_RET_5\ : std_logic ;
  signal \GRLFPC2_0.R.A.AFQ_RET_2\ : std_logic ;
  signal \GRLFPC2_0.R.MK.BUSY_RET\ : std_logic ;
  signal \GRLFPC2_0.R.MK.BUSY_RET_2\ : std_logic ;
  signal \GRLFPC2_0.R.MK.BUSY_RET_3\ : std_logic ;
  signal \GRLFPC2_0.R.MK.BUSY2_RET_1\ : std_logic ;
  signal \GRLFPC2_0.R.A.ST_RET\ : std_logic ;
  signal \GRLFPC2_0.R.A.AFQ_RET_5\ : std_logic ;
  signal \GRLFPC2_0.R.MK.BUSY2_RET\ : std_logic ;
  signal \GRLFPC2_0.R.E.AFSR_RET\ : std_logic ;
  signal \GRLFPC2_0.R.E.SEQERR\ : std_logic ;
  signal \GRLFPC2_0.R.A.SEQERR_RET_3\ : std_logic ;
  signal \GRLFPC2_0.R.A.RS1D\ : std_logic ;
  signal \GRLFPC2_0.R.A.RS2D\ : std_logic ;
  signal \GRLFPC2_0.R.E.AFQ_RET\ : std_logic ;
  signal \GRLFPC2_0.R.I.PC_RET_60\ : std_logic ;
  signal \GRLFPC2_0.R.M.AFSR_RET\ : std_logic ;
  signal \GRLFPC2_0.R.M.AFQ_RET\ : std_logic ;
  signal \GRLFPC2_0.R.E.AFQ_RET_1\ : std_logic ;
  signal \GRLFPC2_0.R.M.AFQ_RET_1\ : std_logic ;
  signal \GRLFPC2_0.R.MK.BUSY2_RET_0_0_A2_0_G0_X\ : std_logic ;
  signal \GRLFPC2_0.R.MK.BUSY_RET_3_0_0_A2_X\ : std_logic ;
  signal \GRLFPC2_0.R.MK.BUSY_RET_2_0_0_A2_0_G0_X\ : std_logic ;
  signal \GRLFPC2_0.R.MK.BUSY2_RET_1_0_0_A2_0_G0\ : std_logic ;
  signal \GRLFPC2_0.R.MK.HOLDN1_0_I_A2_X\ : std_logic ;
  signal \GRLFPC2_0.R.MK.BUSY_RET_4_0_0_A2_0_G0\ : std_logic ;
  signal \GRLFPC2_0.COMB.ANNULFPU_1_U_0_O2\ : std_logic ;
  signal \GRLFPC2_0.COMB.RS1D_1_U\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.FSR.CEXC_1_SN_M3\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.FSR.NONSTD_1_0_X\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN1_FPCI_2_X\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN3_HOLDN_X\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_2_SUM0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW_2_0_65__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD55\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD56\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD57\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_375__G0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_374__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_115__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_58__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SCTRL_NEW_0_0__G0_I_M2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW_6_0_0__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.BUSYMULXFF.UN2_TEMP\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_0_0_13__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW_0_0_7__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW_0_0_7__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_0_0_3__G0_I\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_0_0_2__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_0_0_1__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_76__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_74__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_173__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_243__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_242__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_241__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_240__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_239__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_238__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_237__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_236__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_235__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_234__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_233__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_232__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.STARTSHFT.UN3_NOTRESETORUNIMP\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.STARTSHFT.UN2_NOTDECODEDUNIMP\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN1_TEMP\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN10_S_MOV\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8577_I_0_A2\ : std_logic ;
  signal N_1 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_I_0_0__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.UN36_PCTRL_NEW_I_0_G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_60_SUM0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_60_SUM1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_ADD0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_ADD1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_ADD2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_ADD3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_11\ : std_logic ;
  signal N_30129 : std_logic ;
  signal N_30130 : std_logic ;
  signal N_30132 : std_logic ;
  signal N_30133 : std_logic ;
  signal N_30134 : std_logic ;
  signal N_30135 : std_logic ;
  signal N_30136 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_16\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_18\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_19\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_20\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_21\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_22\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_23\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_24\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_25\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_26\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_27\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_28\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_29\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_30\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_31\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_32\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_33\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_34\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_35\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_36\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_37\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_38\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_39\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_40\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_41\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_42\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_43\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_44\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_45\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_46\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_47\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_48\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_49\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_50\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_51\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_52\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_53\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_54\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_55\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_56\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_11\ : std_logic ;
  signal N_33495_1 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW_6_0_67__G0_I_O4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_47__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_46__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_44__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_41__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_40__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_39__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_35__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_30__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_24__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_23__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_22__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_21__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_20__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_16__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_15__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_14__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_9__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_8__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_2__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_1__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_372__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_319__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_318__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_317__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_316__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_262__G0_I_X4_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_261__G0_I_X4_0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_258__G0_I_X4_0_0_0_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_243__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_242__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_241__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_240__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_239__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_238__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_237__G1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_112__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_111__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_110__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_109__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_108__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_107__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_106__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_105__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_104__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_103__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_102__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_101__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_100__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_99__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_98__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_97__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_96__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_95__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_94__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_93__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_92__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_91__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_90__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_89__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_88__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_87__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_86__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_57__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_55__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_54__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_53__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_52__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_51__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_50__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_49__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_48__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_25__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_24__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_21__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_17__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_16__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_15__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_14__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_13__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_12__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_11__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_10__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_9__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_8__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_7__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_6__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_5__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_4__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_3__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_2__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_1__G2\ : std_logic ;
  signal \GRLFPC2_0.R.I.V_1_0_G2\ : std_logic ;
  signal \GRLFPC2_0.R.I.V_1_0_G0_I_O4\ : std_logic ;
  signal \GRLFPC2_0.R.M.AFQ_RET_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.M.AFSR_RET_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.A.RS2D_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.A.ST_RET_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.E.SEQERR_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.A.RDD_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.A.LD_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.A.FPOP_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.I.EXEC_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.FTT_0_0_2__G1_X\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.FTT_0_0_0__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.NONSTD_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.X.LD_0_0_G1_X\ : std_logic ;
  signal \GRLFPC2_0.R.X.FPOP_0_0_G1_X\ : std_logic ;
  signal \GRLFPC2_0.R.X.AFSR_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.X.AFQ_0_0_G1\ : std_logic ;
  signal \GRLFPC2_0.R.M.LD_0_0_G1_X\ : std_logic ;
  signal \GRLFPC2_0.R.M.FPOP_0_0_G1_X\ : std_logic ;
  signal \GRLFPC2_0.R.E.LD_0_0_G1_X\ : std_logic ;
  signal \GRLFPC2_0.R.E.FPOP_0_0_G1_X\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.RD_0_0_0__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.RD_0_0_1__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.TEM_1_0_0__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.TEM_1_0_1__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.TEM_1_0_2__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.TEM_1_0_3__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.TEM_1_0_4__G1\ : std_logic ;
  signal \GRLFPC2_0.R.STATE_0_0_0__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.FCC_0_0_0__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.FCC_0_0_1__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.CEXC_1_0_0__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.CEXC_1_0_1__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.CEXC_1_0_2__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.CEXC_1_0_3__G1\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.CEXC_1_0_4__G1\ : std_logic ;
  signal \GRLFPC2_0.R.I.CC_0_0_0__G2\ : std_logic ;
  signal \GRLFPC2_0.R.I.CC_0_0_1__G2\ : std_logic ;
  signal \GRLFPC2_0.R.I.EXC_2_0_1__G2\ : std_logic ;
  signal \GRLFPC2_0.R.I.EXC_2_0_2__G2\ : std_logic ;
  signal \GRLFPC2_0.R.I.EXC_2_0_3__G2\ : std_logic ;
  signal \GRLFPC2_0.R.I.EXC_2_0_4__G2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.UN17_U_RDN_I_0_8204_I_A2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.U_RDN_1_8221\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MAPMULXFF.UNIMPMAP_X\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.UN53_SCTRL_NEW\ : std_logic ;
  signal \GRLFPC2_0.N_1213_I_0_O2\ : std_logic ;
  signal \GRLFPC2_0.R.I.RDD_0_0_G1_0_8238_I\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.A.RF1REN_1_8259_I\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.A.RF2REN_1_0_8287_I\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.A.RF2REN_1_8311_I\ : std_logic ;
  signal G_8482 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.TEMP_25\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.TEMP2_0\ : std_logic ;
  signal N_32980_1 : std_logic ;
  signal N_34072_1 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1162\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_9\ : std_logic ;
  signal N_33227_2 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_9_7495\ : std_logic ;
  signal N_33157_1 : std_logic ;
  signal N_28709_1 : std_logic ;
  signal N_29496_1 : std_logic ;
  signal N_34483_1 : std_logic ;
  signal N_28871_1 : std_logic ;
  signal N_34381_1 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8466_I_I_I_X2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11846_I_I_I_X2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_4510_A2_7\ : std_logic ;
  signal NN_1 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_4859_A2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.TOGGLESIG\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.REEXCOVUV.UN20_LOCOV\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXC\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN14_CONDITIONAL\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN30_CONDITIONAL_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SFTLFT.AREGXORBREG_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_8_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_9_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_12_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_11_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.ROMXZSL2FROMC\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_18\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN30_CONDITIONAL_M5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_21\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_24\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPAREGLOADEN_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.A.RF2REN_1_0_8287_I_O4_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN7_RS2V_0_X\ : std_logic ;
  signal \GRLFPC2_0.RS1D_CNST_0_A3_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.RS1_1_SN_M2_I_X\ : std_logic ;
  signal \GRLFPC2_0.RS1D_CNST_0_A2\ : std_logic ;
  signal \GRLFPC2_0.COMB.FPDECODE.RS1D5_0_A2\ : std_logic ;
  signal \GRLFPC2_0.RS1V_0_SQMUXA_1_0_A2_2_X\ : std_logic ;
  signal \GRLFPC2_0.RS1V_0_SQMUXA_1_0_A2_1_X\ : std_logic ;
  signal \GRLFPC2_0.N_939_I_I_2_X\ : std_logic ;
  signal \GRLFPC2_0.COMB.FPDECODE.RS1D5_0_A2_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.RS1V_1_IV\ : std_logic ;
  signal \GRLFPC2_0.RS1V_0_SQMUXA_1_0_A2\ : std_logic ;
  signal \GRLFPC2_0.RS1V_0_SQMUXA_1_0_A2_3_X\ : std_logic ;
  signal \GRLFPC2_0.COMB.FPDECODE.FPOP3_0_A2\ : std_logic ;
  signal \GRLFPC2_0.UN1_FPOP7_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.FPOP_0_0_O2\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.A.RF2REN_1_0_8287_I_A4_0_X\ : std_logic ;
  signal \GRLFPC2_0.N_939_I_I_O2\ : std_logic ;
  signal \GRLFPC2_0.COMB.FPDECODE.FPOP3_0_A2_1_X\ : std_logic ;
  signal \GRLFPC2_0.COMB.FPDECODE.ST_0_A2_0_A2_0_X\ : std_logic ;
  signal \GRLFPC2_0.COMB.RS2D_1_IV_0_O2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_SN_M3_E\ : std_logic ;
  signal NN_2 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19_3_0_.M4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19_3_0_.M3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19_3_0_.M2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN3_NOTAZERODENORM\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN26_NOTBINFNAN\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLAREGEXP.EXPAREGLOADEN_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN1_FPCI_X\ : std_logic ;
  signal \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA_1\ : std_logic ;
  signal \GRLFPC2_0.V.STATE_0_SQMUXA_1_X\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.I.EXEC\ : std_logic ;
  signal \GRLFPC2_0.V.STATE_2_SQMUXA_I_A2_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN1_R.I.V_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN1_MEXC_1\ : std_logic ;
  signal \GRLFPC2_0.R.I.RDD_0_0_G1_0_8238_I_A3\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.STATE\ : std_logic ;
  signal \GRLFPC2_0.UN1_FPCI_21\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.I.EXEC_4_IV_0_A2_X\ : std_logic ;
  signal \GRLFPC2_0.COMB.WREN12_X\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.E.STDATA2_X\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.MK.BUSY_2_4\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_13\ : std_logic ;
  signal \GRLFPC2_0.ANNULRES_0_SQMUXA_10\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN1_FPCI_1_X\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN3_IUEXEC\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.REEXCOVUV.UN3_LOCUV\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CONDMUXMULXFF.UN4_NOTSQRTLFTCC\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.UN3_TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TEMP\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN11_WQSTSETS\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.UN4_TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN4_NOTSHIFTCOUNT1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_SUM0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP_1_C0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.GEN_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP_1_SUM0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN6_NOTPROP_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN10_NOTPROP_0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN27_STKGEN_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_SUM1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN36_STKGEN_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_C1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_C0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN28_STKOUT\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN20_STKOUT\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN22_NOTPROP_0_S\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN16_NOTPROP_0_S\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN18_STKGEN_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.GEN_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.NOTPROP_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_SUM3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN12_STKOUT\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN19_GEN\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN20_GEN\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_C1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.GEN_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_SUM4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_4_M3_E\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_I_M_3950\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_C0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN18_XZXBUS_32_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN18_XZXBUS_40_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN18_XZXBUS_37_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SFTLFT.UN1_GRFPUS\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_AREGSIGN_SEL_INV\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.WQSCTRL_0_3947\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SFTLFT.UN4_TEMP\ : std_logic ;
  signal \GRLFPC2_0.V.STATE_1_SQMUXA_X\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN1_V.STATE\ : std_logic ;
  signal \GRLFPC2_0.COMB.ISFPOP2_1_X\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.FSR.FCC8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLCREGXZ.UN11_INFORCREGSN\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_SUM0\ : std_logic ;
  signal \GRLFPC2_0.COMB.QNE2_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.SEQERR.UN13_OP\ : std_logic ;
  signal \GRLFPC2_0.N_782\ : std_logic ;
  signal \GRLFPC2_0.COMB.SEQERR.SEQERR_0_A3\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.A.AFSR_1_2\ : std_logic ;
  signal \GRLFPC2_0.RS2_0_SQMUXA_3\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN4_LOCK_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.RDD_1.M14_0_O2_0_X\ : std_logic ;
  signal \GRLFPC2_0.COMB.RDD_1.M14_0_A2_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.RDD_1.M14_0_A2_1_X\ : std_logic ;
  signal \GRLFPC2_0.COMB.RDD_1.M14_0_O2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_AREGSIGN_SEL_INV_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DECODESTATUS.UN7_STATUS\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.SELINITREMBIT\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.UN6_U_RDN\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_116_C0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_60_C1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MAPMULXFF.UN4_UNIMPMAP_X\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_2_C0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_58_C0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_114_C0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_10_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.RS2D_1_IV_0_A2_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.RS2D_1_IV_0_O2_0\ : std_logic ;
  signal \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA_X\ : std_logic ;
  signal \GRLFPC2_0.V.FSR.AEXC_1_SQMUXA_X\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN2_INEXACT\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.NOTAM2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN1_S\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN6_S\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.S_CMP\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.STARTSHFT.UN3_NOTDECODEDUNIMP\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.UN17_U_RDN\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN18_XZXBUS_28_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN18_XZXBUS_18_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN18_XZXBUS_19_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN18_XZXBUS_13_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN3_NOTBZERODENORM\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN8_NOTBINFNAN\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN4_NOTAINFNAN\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_60_C0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_114_SUM0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_116_SUM0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_58_SUM0_0\ : std_logic ;
  signal \GRLFPC2_0.WREN1_0_SQMUXA_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_6_M3_E\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.UN132_TEMP_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.UN129_TEMP_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.UN126_TEMP_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.UN120_TEMP_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.UN123_TEMP_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_13_M1_E\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\ : std_logic ;
  signal \GRLFPC2_0.COMB.WREN2_10\ : std_logic ;
  signal \GRLFPC2_0.COMB.WREN1_10_X\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1_0\ : std_logic ;
  signal \GRLFPC2_0.WREN1_1_SQMUXA_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN15_XZROUNDOUT\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLBREGXZ.UN4_XZBREGLOADEN\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN5_SHDVAR\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_8645\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_8715\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_8732\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_8692_TZ\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_9023_TZ\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN7_FEEDBACK_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27_D\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27_D_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_58__G2TT_M2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_58__G2_M9_I_M4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_2_TZ\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_5_TZ\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_5_TZ\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_3_M4_I_X2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_5_TZ\ : std_logic ;
  signal \GRLFPC2_0.COMB.RDD_1.M14_0_A2_2_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.A.RF1REN_1_8259_I_A5_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN1_S_DYADIC_0\ : std_logic ;
  signal \GRLFPC2_0.R.I.V_1_0_G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_2\ : std_logic ;
  signal \GRLFPC2_0.V.FSR.AEXC_1_SQMUXA_0\ : std_logic ;
  signal N_51118 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_2_TZ\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_3_TZ\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_59__G0_XX\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_59__G0_YY\ : std_logic ;
  signal \GRLFPC2_0.COMB.WREN2_9_IV_0\ : std_logic ;
  signal \GRLFPC2_0.UN1_RS1V_0_SQMUXA_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW_6_0_0__G2_0_X\ : std_logic ;
  signal \GRLFPC2_0.RS1V_0_SQMUXA_1_0_A2_2_0\ : std_logic ;
  signal \GRLFPC2_0.RS1D_CNST_0_A2_0\ : std_logic ;
  signal \GRLFPC2_0.RS1D_CNST_0_A3_0_A2_0_0\ : std_logic ;
  signal \GRLFPC2_0.RS1D_CNST_0_A3_0_A2_1_X\ : std_logic ;
  signal \GRLFPC2_0.N_939_I_I_2_0_X\ : std_logic ;
  signal \GRLFPC2_0.COMB.LOCK_1_1_X\ : std_logic ;
  signal \GRLFPC2_0.COMB.RDD_1.M14_0_A2_2_2_X\ : std_logic ;
  signal \GRLFPC2_0.COMB.RDD_1.M14_0_A2_3_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.WREN1_9_IV_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.WREN1_9_IV_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.RDD_1.M14_0_A2_1_0_0_X\ : std_logic ;
  signal \GRLFPC2_0.COMB.RDD_1.M14_0_A2_1_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN8_CCV_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN8_CCV_1\ : std_logic ;
  signal \GRLFPC2_0.RS1V_0_SQMUXA_1_0_A2_0_1\ : std_logic ;
  signal \GRLFPC2_0.RS1V_0_SQMUXA_1_0_A2_0_3\ : std_logic ;
  signal \GRLFPC2_0.R.A.RS2D_0_0_G1_0_X\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G_31_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_11_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN7_FEEDBACK_0_0\ : std_logic ;
  signal \GRLFPC2_0.ANNULRES_0_SQMUXA_10_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN3_IUEXEC_0\ : std_logic ;
  signal \GRLFPC2_0.RS2_0_SQMUXA_2\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN4_LOCK_0_2\ : std_logic ;
  signal \GRLFPC2_0.R.MK.BUSY_RET_4_0_0_A2_0_G0_2\ : std_logic ;
  signal \GRLFPC2_0.V.FSR.FTT_1_SQMUXA_3_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN9_WQSTSETS_0\ : std_logic ;
  signal \GRLFPC2_0.RIN.MK.LDOP_6\ : std_logic ;
  signal \GRLFPC2_0.RIN.MK.LDOP_7\ : std_logic ;
  signal \GRLFPC2_0.RIN.MK.LDOP_8\ : std_logic ;
  signal \GRLFPC2_0.RIN.MK.LDOP_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_3_0\ : std_logic ;
  signal \GRLFPC2_0.N_939_I_I_A2_0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN26_NOTBINFNAN_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN26_NOTBINFNAN_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN26_NOTAINFNAN_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN26_NOTAINFNAN_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN2_INEXACT_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.SEQERR.UN3_QNE_2\ : std_logic ;
  signal \GRLFPC2_0.COMB.SEQERR.UN3_QNE_3\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_13_3\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_13_4\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.MK.RST_1_0_A2_3\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.A.AFQ_1_4\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.A.AFQ_1_6\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.A.AFQ_1_7\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.A.AFQ_1_10\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN1_MEXC_1_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN1_MEXC_1_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN1_FPCI_3_1_X\ : std_logic ;
  signal \GRLFPC2_0.COMB.FPOP_0_0_O2_0_2\ : std_logic ;
  signal \GRLFPC2_0.COMB.ANNULFPU_1_U_0_O2_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.ANNULFPU_1_U_0_O2_1\ : std_logic ;
  signal \GRLFPC2_0.R.I.RDD_0_0_G1_0_8238_I_A3_1\ : std_logic ;
  signal \GRLFPC2_0.R.I.V_1_0_G2_0_0_X\ : std_logic ;
  signal \GRLFPC2_0.R.I.V_1_0_G2_0_3\ : std_logic ;
  signal \GRLFPC2_0.N_939_I_I_A2_1_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_16\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_19\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_20\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_23\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_24\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_27\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_5_M3_E_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_7_M3_E_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_0_X\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_1_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.A.AFSR_1_1_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_3_TZ_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN11_INEXACT_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN12_SRTOSTICKY_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_3_M1_E_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN6_IUEXEC_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_8645_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.A.RF2REN_1_0_8287_I_A4_0_0_X\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.STATE_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.TEMP_25_0\ : std_logic ;
  signal \GRLFPC2_0.N_939_I_I_A2_0_1_X\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.A.RF2REN_1_8311_I_0\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.A.RF1REN_1_8259_I_0\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_0_X\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_14__G2_1\ : std_logic ;
  signal \GRLFPC2_0.R.A.LD_0_0_G1_0\ : std_logic ;
  signal \GRLFPC2_0.R.A.LD_0_0_G1_2_X\ : std_logic ;
  signal \GRLFPC2_0.R.A.LD_0_0_G1_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_44__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLAREGXZ.UN5_XZAREGLOADEN_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_30__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_30__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.ENTRYPOINT_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.ENTRYPOINT_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_23__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_23__G2_2\ : std_logic ;
  signal \GRLFPC2_0.COMB.WREN125_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_5_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_35__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_35__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_16\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_18\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_19\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_22\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_16\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_18\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_21\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_5_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_15__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_15__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_16\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_18\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_19\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_23\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_19\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_19\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_20\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_16\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_18\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_20\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_23\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_24\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_19\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_20\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_21\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_22\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_23\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_18\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_1_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_3_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_16\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_18\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_19\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_39__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_16\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_14\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_16\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_18\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_20\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_22\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_1_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_11\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_10\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_16__G2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_SUM1_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.UN10_U_SNNOTDB_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_9\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_8\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_12\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_13\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_15\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_17\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_19\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_21\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_22\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_23\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_24\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_25\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_27\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_29\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_30\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_31\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_32\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_33\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_35\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_36\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_37\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_38\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_41\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_42\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_45\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_46\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_49\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_50\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_51\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_53\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_55\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN30_CONDITIONAL_M2_E_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN30_CONDITIONAL_M2_E_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1_3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1_5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN30_CONDITIONAL_0_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_0_0_13__G0_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_2_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.BUSYMULXFF.UN2_TEMP_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_4_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_115__G0_0\ : std_logic ;
  signal \GRLFPC2_0.R.I.RDD_0_0_G1_0_8238_I_O4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_C\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\ : std_logic ;
  signal \GRLFPC2_0.WRADDR_1_SQMUXA\ : std_logic ;
  signal \GRLFPC2_0.WRADDR_0_SQMUXA_X\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.FSR.CEXC_1_SN_M2\ : std_logic ;
  signal \GRLFPC2_0.COMB.RDD_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN25_NOTXZYFROMD\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD\ : std_logic ;
  signal \GRLFPC2_0.V.FSR.NONSTD_0_SQMUXA_6_X\ : std_logic ;
  signal \GRLFPC2_0.V.FSR.CEXC_3_SQMUXA\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN1_R.A.RS1_1\ : std_logic ;
  signal \GRLFPC2_0.N_1570_I_I_A2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M11S4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M14S2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5S4\ : std_logic ;
  signal \GRLFPC2_0.COMB.RS1_1_SN_M2_I_A2\ : std_logic ;
  signal \GRLFPC2_0.RS1V_0_SQMUXA_0_A2_X\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G_32\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN1_FPCI_4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_4785_A2_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN6_IUEXEC\ : std_logic ;
  signal G_8368 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPAREGLOADEN\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.FSR.RD_1_SN_M2\ : std_logic ;
  signal \GRLFPC2_0.N_939_I_I_A2\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.A.AFQ_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.V.A.AFSR_1\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN2_HOLDN_0_A2\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR_A\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_7_A\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_A\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN6_IUEXEC_1_A\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_1_A\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_8_A\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN30_CONDITIONAL_M5_A\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_21__G2_A\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_23__G2_2_A\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_6_A\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_7_A\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_13_A\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_17_A\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2_3_A\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_6_A\ : std_logic ;
  signal \GRLFPC2_0.COMB.SEQERR.UN13_OP_A\ : std_logic ;
  signal \GRLFPC2_0.COMB.WREN2_9_IV_0_A\ : std_logic ;
  signal \GRLFPC2_0.COMB.WREN1_9_IV_0_A\ : std_logic ;
  signal \GRLFPC2_0.R.I.V_1_0_G2_0_3_A\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_16_A\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_18_A\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_3_M4_I_X2_A\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_374__G0_A\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.STARTSHFT.UN3_NOTDECODEDUNIMP_A\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1_1_A\ : std_logic ;
  signal \GRLFPC2_0.R.FSR.FTT_0_0_2__G1_A\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_A\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_14_A\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_A\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.GEN_3_A\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_58__G2_M9_I_M4_A\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_0_S\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2_REP1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\ : std_logic ;
  signal \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\ : std_logic ;
  signal \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD_A_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN25_NOTXZYFROMD_RETI\ : std_logic ;
  signal N_10 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_80__G0_A_RETO\ : std_logic ;
  signal N_1_0 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_1_RETO\ : std_logic ;
  signal N_1_1 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO\ : std_logic ;
  signal N_1_2 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_0__G0_0_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_7_RETO\ : std_logic ;
  signal N_1_3 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_78__G0_0_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_2_RETO\ : std_logic ;
  signal N_1_4 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_84__G0_0_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_6_RETO\ : std_logic ;
  signal N_1_5 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_0_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_4_0_RETO\ : std_logic ;
  signal N_1_6 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_6__G0_0_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_1_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\ : std_logic ;
  signal N_1_7 : std_logic ;
  signal N_1_8 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_C_RETO\ : std_logic ;
  signal N_1_9 : std_logic ;
  signal N_1_10 : std_logic ;
  signal N_1_11 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_114__G0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_7\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_6\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_59__G0_XX_MM\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN26_XZYBUSLSBS_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5416_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_2_M1_E_1_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_5_M3_E_1_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_4_M3_E_0_RETI\ : std_logic ;
  signal N_15 : std_logic ;
  signal N_1_12 : std_logic ;
  signal N_1_13 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M11S4_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_A_S_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_6_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5S4_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M2S2_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M8S2_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5S4_1_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M11S4_1_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2_RETI\ : std_logic ;
  signal N_13 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_4_M3_E_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_86__G2_RETO\ : std_logic ;
  signal N_1_14 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_87__G2_RETO\ : std_logic ;
  signal N_1_15 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_88__G2_RETO\ : std_logic ;
  signal N_1_16 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_89__G2_RETO\ : std_logic ;
  signal N_1_17 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_90__G2_RETO\ : std_logic ;
  signal N_1_18 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_91__G2_RETO\ : std_logic ;
  signal N_1_19 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_92__G2_RETO\ : std_logic ;
  signal N_1_20 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_93__G2_RETO\ : std_logic ;
  signal N_1_21 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_94__G2_RETO\ : std_logic ;
  signal N_1_22 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_95__G2_RETO\ : std_logic ;
  signal N_1_23 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_96__G2_RETO\ : std_logic ;
  signal N_1_24 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_97__G2_RETO\ : std_logic ;
  signal N_1_25 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_98__G2_RETO\ : std_logic ;
  signal N_1_26 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_99__G2_RETO\ : std_logic ;
  signal N_1_27 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_100__G2_RETO\ : std_logic ;
  signal N_1_28 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_101__G2_RETO\ : std_logic ;
  signal N_1_29 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_102__G2_RETO\ : std_logic ;
  signal N_1_30 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_103__G2_RETO\ : std_logic ;
  signal N_1_31 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_104__G2_RETO\ : std_logic ;
  signal N_1_32 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_105__G2_RETO\ : std_logic ;
  signal N_1_33 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_106__G2_RETO\ : std_logic ;
  signal N_1_34 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_107__G2_RETO\ : std_logic ;
  signal N_1_35 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_108__G2_RETO\ : std_logic ;
  signal N_1_36 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_109__G2_RETO\ : std_logic ;
  signal N_1_37 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_110__G2_RETO\ : std_logic ;
  signal N_1_38 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_111__G2_RETO\ : std_logic ;
  signal N_1_39 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_112__G2_RETO\ : std_logic ;
  signal N_1_40 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_319__G1_RETO\ : std_logic ;
  signal N_1_41 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_6_M3_E_0_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_7_M3_E_1_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1_RETO\ : std_logic ;
  signal N_1_42 : std_logic ;
  signal N_1_43 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_372__G1_RETO\ : std_logic ;
  signal N_1_44 : std_logic ;
  signal N_14 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN15_XZROUNDOUT_RETI\ : std_logic ;
  signal N_5 : std_logic ;
  signal N_13_0 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_6_M3_E_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_7_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_8_RETI\ : std_logic ;
  signal N_11 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_A_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M14S2_RETI\ : std_logic ;
  signal N_11_0 : std_logic ;
  signal N_12 : std_logic ;
  signal N_11_1 : std_logic ;
  signal N_12_0 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO\ : std_logic ;
  signal N_1_45 : std_logic ;
  signal N_1_46 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_2_0_RETO\ : std_logic ;
  signal N_1_47 : std_logic ;
  signal N_1_48 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_0_RETO\ : std_logic ;
  signal N_1_49 : std_logic ;
  signal N_1_50 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_RETO\ : std_logic ;
  signal N_1_51 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN14_CONDITIONAL_RETO\ : std_logic ;
  signal N_1_52 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_RETO\ : std_logic ;
  signal N_1_53 : std_logic ;
  signal \GRLFPC2_0.R.MK.RST_RET_3\ : std_logic ;
  signal RST_RETO : std_logic ;
  signal N_1_54 : std_logic ;
  signal N_10_0 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_3_M1_E_1_RETI\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_13_M1_E_0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_13_M1_E_RETI\ : std_logic ;
  signal N_16 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_RETO\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT_RETO\ : std_logic ;
  signal N_1_55 : std_logic ;
  signal N_1_56 : std_logic ;
  signal N_2 : std_logic ;
  signal N_3 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_RETI\ : std_logic ;
  signal N_4 : std_logic ;
  signal N_6 : std_logic ;
  signal N_7 : std_logic ;
  signal N_1_57 : std_logic ;
  signal N_1_58 : std_logic ;
  signal N_1_59 : std_logic ;
  signal N_1_60 : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_RETO\ : std_logic ;
  signal N_1_61 : std_logic ;
  signal N_1_62 : std_logic ;
  signal N_1_63 : std_logic ;
  signal N_1_64 : std_logic ;
  signal N_1_65 : std_logic ;
  signal N_1_66 : std_logic ;
  signal N_1_67 : std_logic ;
  signal N_1_68 : std_logic ;
  signal N_1_69 : std_logic ;
  signal N_1_70 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5416\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN26_XZYBUSLSBS\ : std_logic ;
  signal N_1_71 : std_logic ;
  signal N_58149 : std_logic ;
  signal N_58150 : std_logic ;
  signal N_58151 : std_logic ;
  signal N_58152 : std_logic ;
  signal N_58153 : std_logic ;
  signal N_58154 : std_logic ;
  signal N_58155 : std_logic ;
  signal N_58156 : std_logic ;
  signal N_58157 : std_logic ;
  signal N_58158 : std_logic ;
  signal N_58159 : std_logic ;
  signal N_58160 : std_logic ;
  signal N_58161 : std_logic ;
  signal N_58162 : std_logic ;
  signal N_58163 : std_logic ;
  signal N_58164 : std_logic ;
  signal N_58165 : std_logic ;
  signal N_58166 : std_logic ;
  signal N_58167 : std_logic ;
  signal N_58168 : std_logic ;
  signal N_58169 : std_logic ;
  signal N_58170 : std_logic ;
  signal N_58171 : std_logic ;
  signal N_58172 : std_logic ;
  signal N_58173 : std_logic ;
  signal N_58174 : std_logic ;
  signal N_58175 : std_logic ;
  signal N_58176 : std_logic ;
  signal N_58177 : std_logic ;
  signal N_58178 : std_logic ;
  signal N_58179 : std_logic ;
  signal N_58180 : std_logic ;
  signal N_58181 : std_logic ;
  signal N_58182 : std_logic ;
  signal N_58183 : std_logic ;
  signal N_58184 : std_logic ;
  signal N_58185 : std_logic ;
  signal N_58186 : std_logic ;
  signal N_58187 : std_logic ;
  signal N_58188 : std_logic ;
  signal N_58189 : std_logic ;
  signal N_58190 : std_logic ;
  signal N_58191 : std_logic ;
  signal N_58192 : std_logic ;
  signal N_58193 : std_logic ;
  signal N_58194 : std_logic ;
  signal N_58195 : std_logic ;
  signal N_58196 : std_logic ;
  signal N_58197 : std_logic ;
  signal N_58198 : std_logic ;
  signal N_58199 : std_logic ;
  signal N_58200 : std_logic ;
  signal N_58201 : std_logic ;
  signal N_58202 : std_logic ;
  signal N_58203 : std_logic ;
  signal N_58204 : std_logic ;
  signal N_58206 : std_logic ;
  signal N_58207 : std_logic ;
  signal N_58208 : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP2\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_REP0\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_REP1\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_REP2\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_REP3\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_REP4\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_REP5\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP2\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP0\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP1\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\ : std_logic ;
  signal N_58394 : std_logic ;
  signal N_58395 : std_logic ;
  signal N_58396 : std_logic ;
  signal N_58397 : std_logic ;
  signal N_58398 : std_logic ;
  signal N_58399 : std_logic ;
  signal N_58400 : std_logic ;
  signal N_58401 : std_logic ;
  signal N_58402 : std_logic ;
  signal N_58403 : std_logic ;
  signal N_58404 : std_logic ;
  signal N_58405 : std_logic ;
  signal N_58406 : std_logic ;
  signal N_58407 : std_logic ;
  signal N_58408 : std_logic ;
  signal N_58409 : std_logic ;
  signal N_58410 : std_logic ;
  signal N_58411 : std_logic ;
  signal N_58412 : std_logic ;
  signal N_58413 : std_logic ;
  signal N_58414 : std_logic ;
  signal N_58415 : std_logic ;
  signal N_58416 : std_logic ;
  signal N_58417 : std_logic ;
  signal N_58418 : std_logic ;
  signal N_58419 : std_logic ;
  signal N_58420 : std_logic ;
  signal N_58421 : std_logic ;
  signal N_58422 : std_logic ;
  signal N_58423 : std_logic ;
  signal N_58424 : std_logic ;
  signal N_58425 : std_logic ;
  signal N_58426 : std_logic ;
  signal N_58427 : std_logic ;
  signal N_58428 : std_logic ;
  signal N_58429 : std_logic ;
  signal N_58430 : std_logic ;
  signal N_58431 : std_logic ;
  signal N_58432 : std_logic ;
  signal N_58433 : std_logic ;
  signal N_58434 : std_logic ;
  signal N_58435 : std_logic ;
  signal N_58436 : std_logic ;
  signal N_58437 : std_logic ;
  signal N_58438 : std_logic ;
  signal N_58439 : std_logic ;
  signal N_58440 : std_logic ;
  signal N_58441 : std_logic ;
  signal N_58442 : std_logic ;
  signal N_58443 : std_logic ;
  signal N_58444 : std_logic ;
  signal N_58445 : std_logic ;
  signal N_58446 : std_logic ;
  signal N_58447 : std_logic ;
  signal N_58448 : std_logic ;
  signal N_58449 : std_logic ;
  signal N_58450 : std_logic ;
  signal N_58451 : std_logic ;
  signal N_58452 : std_logic ;
  signal N_58453 : std_logic ;
  signal N_58454 : std_logic ;
  signal N_58455 : std_logic ;
  signal N_58456 : std_logic ;
  signal N_58457 : std_logic ;
  signal N_58458 : std_logic ;
  signal N_58459 : std_logic ;
  signal N_58460 : std_logic ;
  signal N_58461 : std_logic ;
  signal N_58462 : std_logic ;
  signal N_58463 : std_logic ;
  signal N_58464 : std_logic ;
  signal N_58465 : std_logic ;
  signal N_58466 : std_logic ;
  signal N_58467 : std_logic ;
  signal N_58468 : std_logic ;
  signal N_58469 : std_logic ;
  signal N_58470 : std_logic ;
  signal N_58471 : std_logic ;
  signal N_58472 : std_logic ;
  signal N_58473 : std_logic ;
  signal N_58474 : std_logic ;
  signal N_58475 : std_logic ;
  signal N_58476 : std_logic ;
  signal N_58477 : std_logic ;
  signal N_58478 : std_logic ;
  signal N_58479 : std_logic ;
  signal N_58480 : std_logic ;
  signal N_58481 : std_logic ;
  signal N_58482 : std_logic ;
  signal N_58483 : std_logic ;
  signal N_58484 : std_logic ;
  signal N_58485 : std_logic ;
  signal N_58486 : std_logic ;
  signal N_58487 : std_logic ;
  signal N_58488 : std_logic ;
  signal N_58489 : std_logic ;
  signal N_58490 : std_logic ;
  signal N_58491 : std_logic ;
  signal N_58492 : std_logic ;
  signal N_58493 : std_logic ;
  signal N_58494 : std_logic ;
  signal N_58495 : std_logic ;
  signal N_58496 : std_logic ;
  signal N_58497 : std_logic ;
  signal N_58498 : std_logic ;
  signal N_58499 : std_logic ;
  signal N_58500 : std_logic ;
  signal N_68349 : std_logic ;
  signal N_68350 : std_logic ;
  signal N_68351 : std_logic ;
  signal HOLDN_INTERNAL : std_logic ;
  signal CPI_DBG_ENABLE_INTERNAL : std_logic ;
  signal CPI_DBG_FSR_INTERNAL : std_logic ;
  signal CPI_DBG_ADDR_INTERNAL : std_logic ;
  signal N_8 : std_logic ;
  signal N_9 : std_logic ;
  signal N_17 : std_logic ;
  signal N_18 : std_logic ;
  signal N_19 : std_logic ;
  signal N_20 : std_logic ;
  signal N_21 : std_logic ;
  signal N_22 : std_logic ;
  signal N_23 : std_logic ;
  signal N_24 : std_logic ;
  signal N_25 : std_logic ;
  signal N_26 : std_logic ;
  signal N_27 : std_logic ;
  signal N_28 : std_logic ;
  signal N_29 : std_logic ;
  signal N_30 : std_logic ;
  signal N_31 : std_logic ;
  signal N_32 : std_logic ;
  signal N_33 : std_logic ;
  signal N_34 : std_logic ;
  signal N_35 : std_logic ;
  signal N_36 : std_logic ;
  signal N_37 : std_logic ;
  signal N_38 : std_logic ;
  signal N_39 : std_logic ;
  signal N_40 : std_logic ;
  signal N_41 : std_logic ;
  signal N_42 : std_logic ;
  signal N_43 : std_logic ;
  signal N_44 : std_logic ;
  signal N_45 : std_logic ;
  signal N_46 : std_logic ;
  signal N_47 : std_logic ;
  signal N_48 : std_logic ;
  signal N_49 : std_logic ;
  signal N_50 : std_logic ;
  signal N_51 : std_logic ;
  signal N_52 : std_logic ;
  signal N_53 : std_logic ;
  signal N_54 : std_logic ;
  signal N_55 : std_logic ;
  signal N_56 : std_logic ;
  signal N_57 : std_logic ;
  signal N_58 : std_logic ;
  signal N_59 : std_logic ;
  signal N_60 : std_logic ;
  signal N_61 : std_logic ;
  signal N_62 : std_logic ;
  signal N_63 : std_logic ;
  signal N_64 : std_logic ;
  signal N_65 : std_logic ;
  signal N_66 : std_logic ;
  signal N_67 : std_logic ;
  signal N_68 : std_logic ;
  signal N_69 : std_logic ;
  signal N_70 : std_logic ;
  signal N_71 : std_logic ;
  signal N_72 : std_logic ;
  signal N_73 : std_logic ;
  signal N_74 : std_logic ;
  signal N_75 : std_logic ;
  signal N_76 : std_logic ;
  signal N_77 : std_logic ;
  signal N_78 : std_logic ;
  signal N_79 : std_logic ;
  signal N_80 : std_logic ;
  signal N_81 : std_logic ;
  signal N_82 : std_logic ;
  signal N_83 : std_logic ;
  signal N_84 : std_logic ;
  signal N_85 : std_logic ;
  signal N_86 : std_logic ;
  signal N_87 : std_logic ;
  signal N_88 : std_logic ;
  signal N_89 : std_logic ;
  signal N_90 : std_logic ;
  signal N_91 : std_logic ;
  signal N_92 : std_logic ;
  signal N_93 : std_logic ;
  signal N_94 : std_logic ;
  signal N_95 : std_logic ;
  signal N_96 : std_logic ;
  signal N_97 : std_logic ;
  signal N_98 : std_logic ;
  signal N_99 : std_logic ;
  signal N_100 : std_logic ;
  signal N_101 : std_logic ;
  signal N_102 : std_logic ;
  signal N_103 : std_logic ;
  signal N_104 : std_logic ;
  signal N_105 : std_logic ;
  signal N_106 : std_logic ;
  signal N_107 : std_logic ;
  signal N_108 : std_logic ;
  signal N_109 : std_logic ;
  signal N_110 : std_logic ;
  signal N_111 : std_logic ;
  signal N_112 : std_logic ;
  signal N_113 : std_logic ;
  signal N_114 : std_logic ;
  signal N_115 : std_logic ;
  signal N_116 : std_logic ;
  signal N_117 : std_logic ;
  signal N_118 : std_logic ;
  signal N_119 : std_logic ;
  signal N_120 : std_logic ;
  signal N_121 : std_logic ;
  signal N_122 : std_logic ;
  signal N_123 : std_logic ;
  signal N_124 : std_logic ;
  signal N_125 : std_logic ;
  signal N_126 : std_logic ;
  signal N_127 : std_logic ;
  signal N_128 : std_logic ;
  signal N_129 : std_logic ;
  signal N_130 : std_logic ;
  signal N_131 : std_logic ;
  signal N_132 : std_logic ;
  signal N_133 : std_logic ;
  signal N_134 : std_logic ;
  signal N_135 : std_logic ;
  signal N_136 : std_logic ;
  signal N_137 : std_logic ;
  signal N_138 : std_logic ;
  signal N_139 : std_logic ;
  signal N_140 : std_logic ;
  signal N_141 : std_logic ;
  signal N_142 : std_logic ;
  signal N_143 : std_logic ;
  signal N_144 : std_logic ;
  signal N_145 : std_logic ;
  signal N_146 : std_logic ;
  signal N_147 : std_logic ;
  signal N_148 : std_logic ;
  signal N_149 : std_logic ;
  signal N_150 : std_logic ;
  signal N_151 : std_logic ;
  signal N_152 : std_logic ;
  signal N_153 : std_logic ;
  signal N_154 : std_logic ;
  signal N_155 : std_logic ;
  signal N_156 : std_logic ;
  signal N_157 : std_logic ;
  signal N_158 : std_logic ;
  signal N_159 : std_logic ;
  signal N_160 : std_logic ;
  signal N_161 : std_logic ;
  signal N_162 : std_logic ;
  signal N_163 : std_logic ;
  signal N_164 : std_logic ;
  signal N_165 : std_logic ;
  signal N_166 : std_logic ;
  signal N_167 : std_logic ;
  signal N_168 : std_logic ;
  signal N_169 : std_logic ;
  signal N_170 : std_logic ;
  signal N_171 : std_logic ;
  signal N_172 : std_logic ;
  signal N_173 : std_logic ;
  signal N_174 : std_logic ;
  signal N_175 : std_logic ;
  signal N_176 : std_logic ;
  signal N_177 : std_logic ;
  signal N_178 : std_logic ;
  signal N_179 : std_logic ;
  signal N_180 : std_logic ;
  signal N_181 : std_logic ;
  signal N_182 : std_logic ;
  signal N_183 : std_logic ;
  signal N_184 : std_logic ;
  signal N_185 : std_logic ;
  signal N_186 : std_logic ;
  signal N_187 : std_logic ;
  signal N_188 : std_logic ;
  signal N_189 : std_logic ;
  signal N_190 : std_logic ;
  signal N_191 : std_logic ;
  signal N_192 : std_logic ;
  signal N_193 : std_logic ;
  signal N_194 : std_logic ;
  signal N_195 : std_logic ;
  signal N_196 : std_logic ;
  signal N_197 : std_logic ;
  signal N_198 : std_logic ;
  signal N_199 : std_logic ;
  signal N_200 : std_logic ;
  signal N_201 : std_logic ;
  signal N_202 : std_logic ;
  signal N_203 : std_logic ;
  signal N_204 : std_logic ;
  signal N_205 : std_logic ;
  signal N_206 : std_logic ;
  signal N_207 : std_logic ;
  signal N_208 : std_logic ;
  signal N_209 : std_logic ;
  signal N_210 : std_logic ;
  signal N_211 : std_logic ;
  signal N_212 : std_logic ;
  signal N_213 : std_logic ;
  signal N_214 : std_logic ;
  signal N_215 : std_logic ;
  signal N_216 : std_logic ;
  signal N_217 : std_logic ;
  signal N_218 : std_logic ;
  signal N_219 : std_logic ;
  signal N_220 : std_logic ;
  signal N_221 : std_logic ;
  signal N_222 : std_logic ;
  signal N_223 : std_logic ;
  signal N_224 : std_logic ;
  signal N_225 : std_logic ;
  signal N_226 : std_logic ;
  signal N_227 : std_logic ;
  signal N_228 : std_logic ;
  signal N_229 : std_logic ;
  signal N_230 : std_logic ;
  signal N_231 : std_logic ;
  signal N_232 : std_logic ;
  signal N_233 : std_logic ;
  signal N_234 : std_logic ;
  signal N_235 : std_logic ;
  signal N_236 : std_logic ;
  signal N_237 : std_logic ;
  signal N_238 : std_logic ;
  signal N_239 : std_logic ;
  signal N_240 : std_logic ;
  signal N_241 : std_logic ;
  signal N_242 : std_logic ;
  signal N_243 : std_logic ;
  signal N_244 : std_logic ;
  signal N_245 : std_logic ;
  signal N_246 : std_logic ;
  signal N_247 : std_logic ;
  signal N_248 : std_logic ;
  signal N_249 : std_logic ;
  signal N_250 : std_logic ;
  signal N_251 : std_logic ;
  signal N_252 : std_logic ;
  signal N_253 : std_logic ;
  signal N_254 : std_logic ;
  signal N_255 : std_logic ;
  signal N_256 : std_logic ;
  signal N_257 : std_logic ;
  signal N_258 : std_logic ;
  signal N_259 : std_logic ;
  signal N_260 : std_logic ;
  signal N_261 : std_logic ;
  signal N_262 : std_logic ;
  signal N_263 : std_logic ;
  signal N_264 : std_logic ;
  signal N_265 : std_logic ;
  signal N_266 : std_logic ;
  signal N_267 : std_logic ;
  signal N_268 : std_logic ;
  signal N_269 : std_logic ;
  signal N_270 : std_logic ;
  signal N_271 : std_logic ;
  signal N_272 : std_logic ;
  signal N_273 : std_logic ;
  signal N_274 : std_logic ;
  signal N_275 : std_logic ;
  signal N_276 : std_logic ;
  signal N_277 : std_logic ;
  signal N_278 : std_logic ;
  signal N_279 : std_logic ;
  signal N_280 : std_logic ;
  signal N_281 : std_logic ;
  signal N_282 : std_logic ;
  signal N_283 : std_logic ;
  signal N_284 : std_logic ;
  signal N_285 : std_logic ;
  signal N_286 : std_logic ;
  signal N_287 : std_logic ;
  signal N_288 : std_logic ;
  signal N_289 : std_logic ;
  signal N_290 : std_logic ;
  signal N_291 : std_logic ;
  signal N_292 : std_logic ;
  signal N_293 : std_logic ;
  signal N_294 : std_logic ;
  signal N_295 : std_logic ;
  signal N_296 : std_logic ;
  signal N_297 : std_logic ;
  signal N_298 : std_logic ;
  signal N_299 : std_logic ;
  signal N_300 : std_logic ;
  signal N_301 : std_logic ;
  signal N_302 : std_logic ;
  signal N_303 : std_logic ;
  signal N_304 : std_logic ;
  signal N_305 : std_logic ;
  signal N_306 : std_logic ;
  signal N_307 : std_logic ;
  signal N_308 : std_logic ;
  signal N_309 : std_logic ;
  signal N_310 : std_logic ;
  signal N_311 : std_logic ;
  signal N_312 : std_logic ;
  signal N_313 : std_logic ;
  signal N_314 : std_logic ;
  signal N_315 : std_logic ;
  signal N_316 : std_logic ;
  signal N_317 : std_logic ;
  signal N_318 : std_logic ;
  signal N_319 : std_logic ;
  signal N_320 : std_logic ;
  signal N_321 : std_logic ;
  signal N_322 : std_logic ;
  signal N_323 : std_logic ;
  signal N_324 : std_logic ;
  signal N_325 : std_logic ;
  signal N_326 : std_logic ;
  signal N_327 : std_logic ;
  signal N_328 : std_logic ;
  signal N_329 : std_logic ;
  signal N_330 : std_logic ;
  signal N_331 : std_logic ;
  signal N_332 : std_logic ;
  signal N_333 : std_logic ;
  signal N_334 : std_logic ;
  signal N_335 : std_logic ;
  signal N_336 : std_logic ;
  signal N_337 : std_logic ;
  signal N_338 : std_logic ;
  signal N_339 : std_logic ;
  signal N_340 : std_logic ;
  signal N_341 : std_logic ;
  signal N_342 : std_logic ;
  signal N_343 : std_logic ;
  signal N_344 : std_logic ;
  signal N_345 : std_logic ;
  signal N_346 : std_logic ;
  signal N_347 : std_logic ;
  signal N_348 : std_logic ;
  signal N_349 : std_logic ;
  signal N_350 : std_logic ;
  signal N_351 : std_logic ;
  signal N_352 : std_logic ;
  signal N_353 : std_logic ;
  signal N_354 : std_logic ;
  signal N_355 : std_logic ;
  signal N_356 : std_logic ;
  signal N_357 : std_logic ;
  signal N_358 : std_logic ;
  signal N_359 : std_logic ;
  signal N_360 : std_logic ;
  signal N_361 : std_logic ;
  signal N_362 : std_logic ;
  signal N_363 : std_logic ;
  signal N_364 : std_logic ;
  signal N_365 : std_logic ;
  signal N_366 : std_logic ;
  signal N_367 : std_logic ;
  signal N_368 : std_logic ;
  signal N_369 : std_logic ;
  signal N_370 : std_logic ;
  signal N_371 : std_logic ;
  signal N_372 : std_logic ;
  signal N_373 : std_logic ;
  signal N_374 : std_logic ;
  signal N_375 : std_logic ;
  signal N_376 : std_logic ;
  signal N_377 : std_logic ;
  signal N_378 : std_logic ;
  signal N_379 : std_logic ;
  signal N_380 : std_logic ;
  signal N_381 : std_logic ;
  signal N_382 : std_logic ;
  signal N_383 : std_logic ;
  signal N_384 : std_logic ;
  signal N_385 : std_logic ;
  signal N_386 : std_logic ;
  signal N_387 : std_logic ;
  signal N_388 : std_logic ;
  signal N_389 : std_logic ;
  signal N_390 : std_logic ;
  signal N_391 : std_logic ;
  signal N_392 : std_logic ;
  signal N_393 : std_logic ;
  signal N_394 : std_logic ;
  signal N_395 : std_logic ;
  signal N_396 : std_logic ;
  signal N_397 : std_logic ;
  signal N_398 : std_logic ;
  signal N_399 : std_logic ;
  signal N_400 : std_logic ;
  signal N_401 : std_logic ;
  signal N_402 : std_logic ;
  signal N_403 : std_logic ;
  signal N_404 : std_logic ;
  signal N_405 : std_logic ;
  signal N_406 : std_logic ;
  signal N_407 : std_logic ;
  signal N_408 : std_logic ;
  signal N_409 : std_logic ;
  signal N_410 : std_logic ;
  signal N_411 : std_logic ;
  signal N_412 : std_logic ;
  signal N_413 : std_logic ;
  signal N_414 : std_logic ;
  signal N_415 : std_logic ;
  signal N_416 : std_logic ;
  signal N_417 : std_logic ;
  signal N_418 : std_logic ;
  signal N_419 : std_logic ;
  signal N_420 : std_logic ;
  signal N_421 : std_logic ;
  signal N_422 : std_logic ;
  signal N_423 : std_logic ;
  signal N_424 : std_logic ;
  signal N_425 : std_logic ;
  signal N_426 : std_logic ;
  signal N_427 : std_logic ;
  signal N_428 : std_logic ;
  signal N_429 : std_logic ;
  signal N_430 : std_logic ;
  signal N_431 : std_logic ;
  signal N_432 : std_logic ;
  signal N_433 : std_logic ;
  signal N_434 : std_logic ;
  signal N_435 : std_logic ;
  signal N_436 : std_logic ;
  signal N_437 : std_logic ;
  signal N_438 : std_logic ;
  signal N_439 : std_logic ;
  signal N_440 : std_logic ;
  signal N_441 : std_logic ;
  signal N_0 : std_logic ;
  signal N_1_72 : std_logic ;
  signal N_2_0 : std_logic ;
  signal N_3_0 : std_logic ;
  signal N_4_0 : std_logic ;
  signal N_5_0 : std_logic ;
  signal N_6_0 : std_logic ;
  signal N_7_0 : std_logic ;
  signal N_8_0 : std_logic ;
  signal N_9_0 : std_logic ;
  signal N_10_1 : std_logic ;
  signal N_11_2 : std_logic ;
  signal N_12_1 : std_logic ;
  signal N_13_1 : std_logic ;
  signal N_14_0 : std_logic ;
  signal N_15_0 : std_logic ;
  signal N_16_0 : std_logic ;
  signal N_17_0 : std_logic ;
  signal N_18_0 : std_logic ;
  signal N_19_0 : std_logic ;
  signal N_20_0 : std_logic ;
  signal N_21_0 : std_logic ;
  signal N_22_0 : std_logic ;
  signal N_23_0 : std_logic ;
  signal N_24_0 : std_logic ;
  signal N_25_0 : std_logic ;
  signal N_26_0 : std_logic ;
  signal N_27_0 : std_logic ;
  signal N_28_0 : std_logic ;
  signal N_29_0 : std_logic ;
  signal N_30_0 : std_logic ;
  signal N_31_0 : std_logic ;
  signal N_32_0 : std_logic ;
  signal N_33_0 : std_logic ;
  signal N_34_0 : std_logic ;
  signal N_35_0 : std_logic ;
  signal N_36_0 : std_logic ;
  signal N_37_0 : std_logic ;
  signal N_38_0 : std_logic ;
  signal N_39_0 : std_logic ;
  signal N_40_0 : std_logic ;
  signal N_41_0 : std_logic ;
  signal N_42_0 : std_logic ;
  signal N_43_0 : std_logic ;
  signal N_44_0 : std_logic ;
  signal N_45_0 : std_logic ;
  signal N_46_0 : std_logic ;
  signal N_47_0 : std_logic ;
  signal N_48_0 : std_logic ;
  signal N_49_0 : std_logic ;
  signal N_50_0 : std_logic ;
  signal N_51_0 : std_logic ;
  signal N_52_0 : std_logic ;
  signal N_53_0 : std_logic ;
  signal N_54_0 : std_logic ;
  signal N_55_0 : std_logic ;
  signal N_56_0 : std_logic ;
  signal N_57_0 : std_logic ;
  signal N_58_0 : std_logic ;
  signal N_59_0 : std_logic ;
  signal N_60_0 : std_logic ;
  signal N_61_0 : std_logic ;
  signal N_62_0 : std_logic ;
  signal N_63_0 : std_logic ;
  signal N_64_0 : std_logic ;
  signal N_65_0 : std_logic ;
  signal N_66_0 : std_logic ;
  signal N_67_0 : std_logic ;
  signal N_68_0 : std_logic ;
  signal N_69_0 : std_logic ;
  signal N_70_0 : std_logic ;
  signal N_71_0 : std_logic ;
  signal N_72_0 : std_logic ;
  signal N_73_0 : std_logic ;
  signal N_74_0 : std_logic ;
  signal N_75_0 : std_logic ;
  signal N_76_0 : std_logic ;
  signal N_77_0 : std_logic ;
  signal N_78_0 : std_logic ;
  signal N_79_0 : std_logic ;
  signal N_80_0 : std_logic ;
  signal N_81_0 : std_logic ;
  signal N_82_0 : std_logic ;
  signal N_83_0 : std_logic ;
  signal N_84_0 : std_logic ;
  signal N_85_0 : std_logic ;
  signal N_86_0 : std_logic ;
  signal N_87_0 : std_logic ;
  signal N_88_0 : std_logic ;
  signal N_89_0 : std_logic ;
  signal N_90_0 : std_logic ;
  signal N_91_0 : std_logic ;
  signal N_92_0 : std_logic ;
  signal N_93_0 : std_logic ;
  signal N_94_0 : std_logic ;
  signal N_95_0 : std_logic ;
  signal N_96_0 : std_logic ;
  signal N_97_0 : std_logic ;
  signal N_98_0 : std_logic ;
  signal N_99_0 : std_logic ;
  signal N_100_0 : std_logic ;
  signal N_101_0 : std_logic ;
  signal N_102_0 : std_logic ;
  signal N_103_0 : std_logic ;
  signal N_104_0 : std_logic ;
  signal N_105_0 : std_logic ;
  signal N_106_0 : std_logic ;
  signal N_107_0 : std_logic ;
  signal N_108_0 : std_logic ;
  signal N_109_0 : std_logic ;
  signal N_110_0 : std_logic ;
  signal N_111_0 : std_logic ;
  signal N_112_0 : std_logic ;
  signal N_113_0 : std_logic ;
  signal N_114_0 : std_logic ;
  signal N_115_0 : std_logic ;
  signal N_116_0 : std_logic ;
  signal N_117_0 : std_logic ;
  signal N_118_0 : std_logic ;
  signal N_119_0 : std_logic ;
  signal N_120_0 : std_logic ;
  signal N_121_0 : std_logic ;
  signal N_122_0 : std_logic ;
  signal N_123_0 : std_logic ;
  signal N_124_0 : std_logic ;
  signal N_125_0 : std_logic ;
  signal N_126_0 : std_logic ;
  signal N_127_0 : std_logic ;
  signal N_128_0 : std_logic ;
  signal N_129_0 : std_logic ;
  signal N_130_0 : std_logic ;
  signal N_131_0 : std_logic ;
  signal N_132_0 : std_logic ;
  signal N_133_0 : std_logic ;
  signal N_134_0 : std_logic ;
  signal N_135_0 : std_logic ;
  signal N_136_0 : std_logic ;
  signal N_137_0 : std_logic ;
  signal N_138_0 : std_logic ;
  signal N_139_0 : std_logic ;
  signal N_140_0 : std_logic ;
  signal N_141_0 : std_logic ;
  signal N_142_0 : std_logic ;
  signal N_143_0 : std_logic ;
  signal N_144_0 : std_logic ;
  signal N_145_0 : std_logic ;
  signal N_146_0 : std_logic ;
  signal N_147_0 : std_logic ;
  signal N_148_0 : std_logic ;
  signal N_149_0 : std_logic ;
  signal N_150_0 : std_logic ;
  signal N_151_0 : std_logic ;
  signal N_152_0 : std_logic ;
  signal N_153_0 : std_logic ;
  signal N_154_0 : std_logic ;
  signal N_155_0 : std_logic ;
  signal N_156_0 : std_logic ;
  signal N_157_0 : std_logic ;
  signal N_158_0 : std_logic ;
  signal N_159_0 : std_logic ;
  signal N_160_0 : std_logic ;
  signal N_161_0 : std_logic ;
  signal N_162_0 : std_logic ;
  signal N_163_0 : std_logic ;
  signal N_606 : std_logic ;
  signal N_607 : std_logic ;
  signal N_608 : std_logic ;
  signal N_609 : std_logic ;
  signal N_610 : std_logic ;
  signal N_611 : std_logic ;
  signal N_612 : std_logic ;
  signal N_613 : std_logic ;
  signal N_614 : std_logic ;
  signal N_615 : std_logic ;
  signal N_616 : std_logic ;
  signal N_617 : std_logic ;
  signal N_618 : std_logic ;
  signal N_619 : std_logic ;
  signal N_620 : std_logic ;
  signal N_621 : std_logic ;
  signal N_622 : std_logic ;
  signal N_623 : std_logic ;
  signal N_624 : std_logic ;
  signal N_625 : std_logic ;
  signal N_626 : std_logic ;
  signal N_627 : std_logic ;
  signal N_628 : std_logic ;
  signal N_629 : std_logic ;
  signal N_630 : std_logic ;
  signal N_631 : std_logic ;
  signal N_632 : std_logic ;
  signal N_633 : std_logic ;
  signal N_634 : std_logic ;
  signal N_635 : std_logic ;
  signal N_636 : std_logic ;
  signal N_637 : std_logic ;
  signal N_638 : std_logic ;
  signal N_639 : std_logic ;
  signal N_640 : std_logic ;
  signal N_641 : std_logic ;
  signal N_642 : std_logic ;
  signal N_643 : std_logic ;
  signal N_644 : std_logic ;
  signal N_645 : std_logic ;
  signal N_646 : std_logic ;
  signal N_647 : std_logic ;
  signal N_648 : std_logic ;
  signal N_649 : std_logic ;
  signal N_650 : std_logic ;
  signal N_651 : std_logic ;
  signal N_652 : std_logic ;
  signal N_653 : std_logic ;
  signal N_654 : std_logic ;
  signal N_655 : std_logic ;
  signal N_656 : std_logic ;
  signal N_657 : std_logic ;
  signal N_658 : std_logic ;
  signal N_659 : std_logic ;
  signal N_660 : std_logic ;
  signal N_661 : std_logic ;
  signal N_662 : std_logic ;
  signal N_663 : std_logic ;
  signal N_664 : std_logic ;
  signal N_665 : std_logic ;
  signal N_666 : std_logic ;
  signal N_667 : std_logic ;
  signal N_668 : std_logic ;
  signal N_669 : std_logic ;
  signal N_670 : std_logic ;
  signal N_671 : std_logic ;
  signal N_672 : std_logic ;
  signal N_673 : std_logic ;
  signal N_674 : std_logic ;
  signal N_675 : std_logic ;
  signal N_676 : std_logic ;
  signal N_677 : std_logic ;
  signal N_678 : std_logic ;
  signal N_679 : std_logic ;
  signal N_680 : std_logic ;
  signal N_681 : std_logic ;
  signal N_682 : std_logic ;
  signal N_683 : std_logic ;
  signal N_684 : std_logic ;
  signal N_685 : std_logic ;
  signal N_686 : std_logic ;
  signal N_687 : std_logic ;
  signal N_688 : std_logic ;
  signal N_689 : std_logic ;
  signal N_690 : std_logic ;
  signal N_691 : std_logic ;
  signal N_692 : std_logic ;
  signal N_693 : std_logic ;
  signal N_694 : std_logic ;
  signal N_695 : std_logic ;
  signal N_696 : std_logic ;
  signal N_697 : std_logic ;
  signal N_698 : std_logic ;
  signal N_699 : std_logic ;
  signal N_700 : std_logic ;
  signal N_701 : std_logic ;
  signal N_702 : std_logic ;
  signal N_703 : std_logic ;
  signal N_704 : std_logic ;
  signal N_705 : std_logic ;
  signal N_706 : std_logic ;
  signal N_707 : std_logic ;
  signal N_708 : std_logic ;
  signal N_709 : std_logic ;
  signal N_710 : std_logic ;
  signal N_711 : std_logic ;
  signal N_712 : std_logic ;
  signal N_713 : std_logic ;
  signal N_714 : std_logic ;
  signal N_715 : std_logic ;
  signal N_716 : std_logic ;
  signal N_717 : std_logic ;
  signal N_718 : std_logic ;
  signal N_719 : std_logic ;
  signal N_720 : std_logic ;
  signal N_721 : std_logic ;
  signal N_722 : std_logic ;
  signal N_723 : std_logic ;
  signal N_724 : std_logic ;
  signal N_725 : std_logic ;
  signal N_726 : std_logic ;
  signal N_727 : std_logic ;
  signal N_728 : std_logic ;
  signal N_729 : std_logic ;
  signal N_730 : std_logic ;
  signal N_731 : std_logic ;
  signal N_732 : std_logic ;
  signal N_733 : std_logic ;
  signal \GRLFPC2_0.COMB.V.A.AFQ_1_I\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\ : std_logic ;
  signal \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\ : std_logic ;
  signal \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\ : std_logic ;
  signal \GRLFPC2_0.FPI.LDOP_I\ : std_logic ;
  signal CPO_EXCZ : std_logic ;
  signal CPO_CCVZ : std_logic ;
  signal CPO_LDLOCKZ : std_logic ;
  signal CPO_HOLDNZ : std_logic ;
  signal RFI1_REN1Z : std_logic ;
  signal RFI1_REN2Z : std_logic ;
  signal RFI1_WRENZ : std_logic ;
  signal RFI2_REN1Z : std_logic ;
  signal RFI2_REN2Z : std_logic ;
  signal RFI2_WRENZ : std_logic ;
begin
VCC <= '1';
GND <= '0';
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIU736_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58500,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_1_RNI31EU3_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(110),
cin => N_58499);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIV736_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58498,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_3_RNI0O5O3_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(109),
cin => N_58497);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNI7PE2_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58496,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_3_RNITVDH3_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(108),
cin => N_58495);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNI8TE2_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58494,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_1_RNINFAL3_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(107),
cin => N_58493);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNI91F2_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58492,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(12));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_3_RNIKO8H4_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(106),
cin => N_58491);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIA5F2_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58490,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(13));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_3_RNIFUB16_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(105),
cin => N_58489);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIB9F2_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58488,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(14));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_2_RNIGJC67_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(104),
cin => N_58487);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNICDF2_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58486,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(15));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_3_RNIRECF7_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(103),
cin => N_58485);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIDHF2_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58484,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(16));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_1_RNIUTVU6_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(102),
cin => N_58483);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIELF2_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58482,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(17));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_3_RNI1EKR5_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(101),
cin => N_58481);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNI8PE2_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58480,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(20));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_2_RNIOKSC4_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(98),
cin => N_58479);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNI9TE2_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58478,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(21));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_3_RNIP8L54_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(97),
cin => N_58477);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIA1F2_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58476,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(22));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_2_RNI2SU54_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(96),
cin => N_58475);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIB5F2_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58474,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(23));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_1_RNI90JT3_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(95),
cin => N_58473);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIC9F2_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58472,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(24));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_3_RNI09K04_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(94),
cin => N_58471);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIDDF2_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58470,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(25));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_2_RNIRDGB4_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(93),
cin => N_58469);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIEHF2_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58468,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(26));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_3_RNID7VQ4_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(92),
cin => N_58467);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIFLF2_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58466,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(27));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_2_RNI8LT55_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(91),
cin => N_58465);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIGPF2_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58464,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(28));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_3_RNITV545_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(90),
cin => N_58463);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIHTF2_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58462,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(29));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_RNILEET4_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(89),
cin => N_58461);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNI9PE2_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58460,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(30));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_RNIPDME4_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(88),
cin => N_58459);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIATE2_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58458,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(31));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_1_RNIMVN84_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(87),
cin => N_58457);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIB1F2_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58456,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(32));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_1_RNIRGA84_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(86),
cin => N_58455);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIS736_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58454,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_2_RNIHG744_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(112),
cin => N_58453);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIT736_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58452,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(7));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_1_RNIPUJ24_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(111),
cin => N_58451);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIEDF2_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58450,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(35));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_3_RNIH7GC4_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(83),
cin => N_58449);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIFHF2_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58448,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(36));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_RNIGOBC4_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(82),
cin => N_58447);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIGLF2_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58446,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(37));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_2_RNIC27E4_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(81),
cin => N_58445);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIHPF2_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58444,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(38));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_1_RNI9BK14_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(80),
cin => N_58443);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIITF2_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58442,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(39));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_RNI003R3_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(79),
cin => N_58441);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIAPE2_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58440,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(40));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_1_RNII8I04_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(78),
cin => N_58439);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIBTE2_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58438,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(41));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_RNIUG6O3_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(77),
cin => N_58437);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIC1F2_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58436,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(42));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_2_RNIB65I3_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(76),
cin => N_58435);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNID5F2_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58434,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(43));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_RNIVTRD3_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(75),
cin => N_58433);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIE9F2_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58432,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(44));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_2_RNICN8K3_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(74),
cin => N_58431);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIFDF2_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58430,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(45));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_2_RNIF0JT3_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(73),
cin => N_58429);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIGHF2_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58428,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(46));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_3_RNIC4G04_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(72),
cin => N_58427);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIHLF2_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58426,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(47));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_3_RNIBD014_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(71),
cin => N_58425);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIFPF2_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58424,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(18));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_1_RNI2KVP4_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(100),
cin => N_58423);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIGTF2_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58422,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(19));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_RNI4CDF4_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(99),
cin => N_58421);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIIPF2_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58420,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(48));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_1_RNI0FT64_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(70),
cin => N_58419);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIJTF2_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58418,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(49));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_1_RNIMG654_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(69),
cin => N_58417);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIBPE2_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58416,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(50));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_3_RNI9N4O3_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(68),
cin => N_58415);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNICTE2_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58414,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(51));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_RNI77NC3_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(67),
cin => N_58413);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNID1F2_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58412,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(52));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_3_RNIT93F3_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(66),
cin => N_58411);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIE5F2_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58410,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(53));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_3_RNIGKEF3_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(65),
cin => N_58409);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIF9F2_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58408,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(54));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_RNI7CCO3_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(64),
cin => N_58407);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIGDF2_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58406,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(55));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_2_RNI7CTR3_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(63),
cin => N_58405);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIHHF2_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58404,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(56));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_3_RNI345R3_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(62),
cin => N_58403);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIILF2_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58402,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(57));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_3_RNIVFBG3_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(61),
cin => N_58401);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIC5F2_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58400,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(33));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_1_RNI7NR24_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(85),
cin => N_58399);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNID9F2_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58398,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(34));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_3_RNID2884_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(84),
cin => N_58397);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_ADD0_START: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58396,
dataa => VCC);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD0_START: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58395,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN8_TEMP_U\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_ADD0_START: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_58394,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.MIXOIN\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_26_RNIB63E1_7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_6__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_26_RNIB63E1_4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_6__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_26_RNIB63E1_5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_6__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_26_RNIB63E1_6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_6__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_26_RNIB63E1_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_6__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_26_RNIB63E1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_6__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_26_RNIB63E1_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_6__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_26_RNIB63E1_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_6__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_14_RNI663E1_7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_7_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_0__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_14_RNI663E1_5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_7_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_0__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_14_RNI663E1_6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_7_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_0__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_14_RNI663E1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_7_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_0__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_14_RNI663E1_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_7_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_0__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_14_RNI663E1_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_7_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_0__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_14_RNI663E1_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_7_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_0__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_14_RNI663E1_4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_7_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_0__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_20_RNI70DC1_5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_U_RETO\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_6_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_84__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_20_RNI70DC1_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_U_RETO\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_6_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_84__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_20_RNI70DC1_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_U_RETO\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_6_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_84__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_20_RNI70DC1_7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_U_RETO\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_6_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_84__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_20_RNI70DC1_4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_U_RETO\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_6_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_84__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_20_RNI70DC1_6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_U_RETO\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_6_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_84__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_20_RNI70DC1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_U_RETO\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_6_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_84__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_20_RNI70DC1_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_U_RETO\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_6_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_84__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_8_RNIR9B12_7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_RETO\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_C_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_1_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_8_RNIR9B12_6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_RETO\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_C_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_1_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_8_RNIR9B12: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_RETO\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_C_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_1_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_8_RNIR9B12_4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_RETO\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_C_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_1_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_8_RNIR9B12_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_RETO\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_C_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_1_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_8_RNIR9B12_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_RETO\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_C_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_1_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_8_RNIR9B12_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_RETO\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_C_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_1_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_8_RNIR9B12_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_RETO\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_C_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_1_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_12_RNIPRP02_5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_M_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_12_RNIPRP02_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_M_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_12_RNIPRP02_6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_M_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_12_RNIPRP02_4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_M_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_12_RNIPRP02_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_M_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_12_RNIPRP02_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_M_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_12_RNIPRP02_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_M_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_23_RNI463E1_4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_4_0_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_23_RNI463E1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_4_0_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_23_RNI463E1_6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_4_0_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_23_RNI463E1_5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_4_0_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_23_RNI463E1_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_4_0_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_23_RNI463E1_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_4_0_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_23_RNI463E1_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_4_0_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_23_RNI463E1_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_4_0_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_4_RNIN52O1_7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_X_RETO\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_80__G0_A_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_4_RNIN52O1_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_X_RETO\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_80__G0_A_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_4_RNIN52O1_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_X_RETO\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_80__G0_A_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_4_RNIN52O1_5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_X_RETO\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_80__G0_A_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_4_RNIN52O1_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_X_RETO\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_80__G0_A_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_4_RNIN52O1_6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_X_RETO\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_80__G0_A_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_4_RNIN52O1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_X_RETO\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_80__G0_A_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_4_RNIN52O1_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_X_RETO\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_80__G0_A_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_17_RNIT0DC1_5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_2_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_78__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_17_RNIT0DC1_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_2_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_78__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_17_RNIT0DC1_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_2_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_78__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_17_RNIT0DC1_4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_2_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_78__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_17_RNIT0DC1_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_2_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_78__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_17_RNIT0DC1_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_2_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_78__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_17_RNIT0DC1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_2_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_78__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_17_RNII63E1_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_2_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_78__G0_0_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIGOP2_1_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(5),
datab => \GRLFPC2_0.FPI.LDOP_REP5\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIGOP2_0_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(5),
datab => \GRLFPC2_0.FPI.LDOP_REP5\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_REP2_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010011000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_REP1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010011000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_REP2_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010011000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_REP1_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010011000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_116_REP1_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_REP2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP2\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_REP1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_118_REP2_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP2\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_118_REP1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP1\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN50_ZERO_REP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111001111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN50_ZERO_REP1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111001111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_0_REP1_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011110111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN20_ZERO_REP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111001111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN20_ZERO_REP1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111001111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_0_REP1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010111001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN35_ZERO_REP1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111001111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_0_REP1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010111001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN5_ZERO_REP1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_A\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_REP2_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111101000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(43),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_REP1_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111101000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(43),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_RNIGPS6_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TEMP\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD10\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD11\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN12_SRTOSTICKY_3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIJE8B_0_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_REP1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLAREGXZ.UN5_XZAREGLOADEN_0\,
datac => \GRLFPC2_0.FPI.LDOP_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.WQSCTRL_0\(67));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_REP0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLAREGXZ.UN5_XZAREGLOADEN_0\,
datac => \GRLFPC2_0.FPI.LDOP_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.WQSCTRL_0\(67));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_REP4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN1_TEMP\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW\(77),
datad => \GRLFPC2_0.FPI.LDOP_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_REP3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN1_TEMP\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW\(77),
datad => \GRLFPC2_0.FPI.LDOP_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_REP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN1_TEMP\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW\(77),
datad => \GRLFPC2_0.FPI.LDOP_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_REP1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN1_TEMP\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW\(77),
datad => \GRLFPC2_0.FPI.LDOP_REP1\);
GRLFPC2_0_FPI_LDOP_REP5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.FPI.LDOP_REP5\,
dataa => \GRLFPC2_0.RIN.MK.LDOP_7\,
datab => \GRLFPC2_0.RIN.MK.LDOP_8\,
datac => \GRLFPC2_0.RIN.MK.LDOP_9\,
datad => \GRLFPC2_0.FPI.LDOP_0_X\);
GRLFPC2_0_FPI_LDOP_REP4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.FPI.LDOP_REP4\,
dataa => \GRLFPC2_0.RIN.MK.LDOP_7\,
datab => \GRLFPC2_0.RIN.MK.LDOP_8\,
datac => \GRLFPC2_0.RIN.MK.LDOP_9\,
datad => \GRLFPC2_0.FPI.LDOP_0_X\);
GRLFPC2_0_FPI_LDOP_REP3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.FPI.LDOP_REP3\,
dataa => \GRLFPC2_0.RIN.MK.LDOP_7\,
datab => \GRLFPC2_0.RIN.MK.LDOP_8\,
datac => \GRLFPC2_0.RIN.MK.LDOP_9\,
datad => \GRLFPC2_0.FPI.LDOP_0_X\);
GRLFPC2_0_FPI_LDOP_REP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.FPI.LDOP_REP2\,
dataa => \GRLFPC2_0.RIN.MK.LDOP_7\,
datab => \GRLFPC2_0.RIN.MK.LDOP_8\,
datac => \GRLFPC2_0.RIN.MK.LDOP_9\,
datad => \GRLFPC2_0.FPI.LDOP_0_X\);
GRLFPC2_0_FPI_LDOP_REP1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.FPI.LDOP_REP1\,
dataa => \GRLFPC2_0.RIN.MK.LDOP_7\,
datab => \GRLFPC2_0.RIN.MK.LDOP_8\,
datac => \GRLFPC2_0.RIN.MK.LDOP_9\,
datad => \GRLFPC2_0.FPI.LDOP_0_X\);
GRLFPC2_0_FPI_LDOP_REP0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.FPI.LDOP_REP0\,
dataa => \GRLFPC2_0.RIN.MK.LDOP_7\,
datab => \GRLFPC2_0.RIN.MK.LDOP_8\,
datac => \GRLFPC2_0.RIN.MK.LDOP_9\,
datad => \GRLFPC2_0.FPI.LDOP_0_X\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIN7RL_1_71_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011111101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(72),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(71),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIN7RL_0_71_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011111101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(72),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(71),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN38_SHDVAR_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5416_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_57__G2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA_0_RNI33PF: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_115__G0_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_0\,
datac => \GRLFPC2_0.FPI.LDOP_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN15_XZROUNDOUT: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN15_XZROUNDOUT_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_0_0_3__G0_I\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPYBUS_2_1_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2_1_RETI\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW\(10),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_30__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_249_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(249),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(60),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\(249),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_246_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(246),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\(246),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_248_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(248),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\(248),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_247_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(247),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\(247),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_245_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(245),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(245),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\(245),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_5_RNINQ4I: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
dataa => \GRLFPC2_0.FPI.LDOP_RETO\,
datab => RFO2_DATA1_RETO(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(85));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_3_RNIKQ4I: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
dataa => \GRLFPC2_0.FPI.LDOP_RETO\,
datab => RFO2_DATA1_RETO(28),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(84));
\GRLFPC2_0_R_FSR_TEM_RNO_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.R.FSR.TEM_1_0_0__G1\,
dataa => N_8,
datab => N_433,
datac => \GRLFPC2_0.COMB.V.FSR.RD_1_SN_M2\,
datad => \GRLFPC2_0.COMB.V.FSR.TEM_1_0_X\(0));
\GRLFPC2_0_R_FSR_RD_RNO_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.R.FSR.RD_0_0_0__G1\,
dataa => N_8,
datab => N_440,
datac => \GRLFPC2_0.COMB.V.FSR.RD_1_SN_M2\,
datad => \GRLFPC2_0.COMB.V.FSR.RD_1_0_X\(0));
GRLFPC2_0_R_FSR_NONSTD_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.R.FSR.NONSTD_0_0_G1\,
dataa => N_8,
datab => N_432,
datac => \GRLFPC2_0.COMB.V.FSR.RD_1_SN_M2\,
datad => \GRLFPC2_0.COMB.V.FSR.NONSTD_1_0_X\);
\GRLFPC2_0_R_FSR_TEM_RNO_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.R.FSR.TEM_1_0_2__G1\,
dataa => N_8,
datab => N_435,
datac => \GRLFPC2_0.COMB.V.FSR.RD_1_SN_M2\,
datad => \GRLFPC2_0.COMB.V.FSR.TEM_1_0_X\(2));
\GRLFPC2_0_R_FSR_TEM_RNO_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.R.FSR.TEM_1_0_3__G1\,
dataa => N_8,
datab => N_436,
datac => \GRLFPC2_0.COMB.V.FSR.RD_1_SN_M2\,
datad => \GRLFPC2_0.COMB.V.FSR.TEM_1_0_X\(3));
\GRLFPC2_0_R_FSR_TEM_RNO_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.R.FSR.TEM_1_0_4__G1\,
dataa => N_8,
datab => N_437,
datac => \GRLFPC2_0.COMB.V.FSR.RD_1_SN_M2\,
datad => \GRLFPC2_0.COMB.V.FSR.TEM_1_0_X\(4));
\GRLFPC2_0_R_FSR_TEM_RNO_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.R.FSR.TEM_1_0_1__G1\,
dataa => N_8,
datab => N_434,
datac => \GRLFPC2_0.COMB.V.FSR.RD_1_SN_M2\,
datad => \GRLFPC2_0.COMB.V.FSR.TEM_1_0_X\(1));
\GRLFPC2_0_R_FSR_RD_RNO_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.R.FSR.RD_0_0_1__G1\,
dataa => N_8,
datab => N_441,
datac => \GRLFPC2_0.COMB.V.FSR.RD_1_SN_M2\,
datad => \GRLFPC2_0.COMB.V.FSR.RD_1_0_X\(1));
RETGRLFPC2_0_COMB_ANNULFPU_1_U_0_O2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110100")
port map (
combout => N_58208,
dataa => \GRLFPC2_0.COMB.UN1_FPCI_X\,
datab => \GRLFPC2_0.R.X.SEQERR\,
datac => \GRLFPC2_0.COMB.ANNULFPU_1_U_0_O2_1\,
datad => \GRLFPC2_0.COMB.ANNULFPU_1_U_0_O2_0\);
RETGRLFPC2_0_COMB_V_MK_RST_1_0_A2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => N_58207,
dataa => \GRLFPC2_0.R.MK.HOLDN2\,
datab => \GRLFPC2_0.R.MK.RST_RET_6\,
datac => \GRLFPC2_0.R.MK.RST2\,
datad => \GRLFPC2_0.COMB.V.MK.RST_1_0_A2_3\);
RETGRLFPC2_0_N_939_I_I_A2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => N_58206,
dataa => N_89,
datab => N_90,
datac => \GRLFPC2_0.N_939_I_I_A2_0_1_X\,
datad => \GRLFPC2_0.N_939_I_I_O2\);
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23_1_SUM_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011101111000")
port map (
combout => N_58204,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_114_C0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_0\(56));
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_0_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100111110101111")
port map (
combout => N_58203,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.UN10_U_SNNOTDB_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.TOGGLESIG\);
RETGRLFPC2_0_FPI_LDOP_0_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110111111101")
port map (
combout => N_58202,
dataa => N_8,
datab => \GRLFPC2_0.R.MK.RST2\,
datac => \GRLFPC2_0.COMB.V.MK.RST_1_0_A2\);
RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_UN10_SELECTEDMIPTR: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => N_58201,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CONDMUXMULXFF.UN4_NOTSQRTLFTCC\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27\);
RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_D: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001111110001")
port map (
combout => N_58200,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CONDMUXMULXFF.UN4_NOTSQRTLFTCC\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27\);
RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_C: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110011001100")
port map (
combout => N_58199,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.UN4_TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.TEMP_25\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.STARTSHFT.UN3_NOTRESETORUNIMP\);
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => N_58198,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2\);
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M_0_57__G2\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => N_58197,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(57));
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M_0_56__G2\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => N_58196,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(56));
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => N_58195,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_55__G2\);
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => N_58194,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_25__G2\);
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_58__G0\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010101000000")
port map (
combout => N_58193,
dataa => \GRLFPC2_0.FPI.LDOP_REP5\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_317__G1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_58__G2_M9_I_M4\);
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => N_58192,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1\(11));
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => N_58191,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_8__G2\);
RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN16_NOTXZYFROMD_REP1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => N_58190,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(1));
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_0_84__G0_I_A3\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111011101110111")
port map (
combout => N_58189,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.LDOP_REP5\);
RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => N_58188,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_0\,
datac => \GRLFPC2_0.FPI.LDOP_REP5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP1\);
RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA_REP1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => N_58187,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_0\,
datac => \GRLFPC2_0.FPI.LDOP_REP5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP1\);
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_372__G1\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100110001001100")
port map (
combout => N_58186,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP2\(2));
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => N_58185,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_54__G2\);
RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_SN_M4_0_REP1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100110010")
port map (
combout => N_58184,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1_RETI\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN25_NOTXZYFROMD_RETI\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1_RETI\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD_RETI\);
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M_0_2__G2\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => N_58183,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(2));
RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M11S4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => N_58182,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_4__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_3__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_5__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_6__G2\);
RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M5S4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => N_58181,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_14__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_11__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_12__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_13__G2\);
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O19_2_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110111011101")
port map (
combout => N_58180,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83));
RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110111111101")
port map (
combout => N_58179,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CONDMUXMULXFF.UN4_NOTSQRTLFTCC\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27\);
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_0_84__G0\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => N_58178,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_U_RETO\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_6_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_84__G0_0_RETO\);
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_7_1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => N_58177,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84));
RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN14_CONDITIONAL: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111000000000")
port map (
combout => N_58176,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_4\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_5\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN3_NOTAZERODENORM\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS\(3));
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000010101")
port map (
combout => N_58175,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN3_NOTBZERODENORM\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN26_NOTBINFNAN\);
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => N_58174,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_4\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_5\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN3_NOTBZERODENORM\);
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_IV_I_0_6__G0\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => N_58173,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_6__G0_0_RETO\);
RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN53_SCTRL_NEW: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000110101")
port map (
combout => N_58172,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.U_RDN_1\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW\(9));
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_REP1EN_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => N_58171,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_16__G2\);
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => N_58170,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_16__G2\);
RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN15_NOTXZYFROMD_0_REP1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110010100000")
port map (
combout => N_58169,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_375__G0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(11));
RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN25_NOTXZYFROMD: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010001000")
port map (
combout => N_58168,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_374__G0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(12),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(11));
RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN15_NOTXZYFROMD: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011110010")
port map (
combout => N_58167,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1_RETI\);
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_115__G0\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000010001000")
port map (
combout => N_58166,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_115__G0_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(115),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(115),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => N_58165,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2\);
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100011001000")
port map (
combout => N_58164,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.UN53_SCTRL_NEW\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1I\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_0_0_3__G0_I\);
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => N_58163,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_52__G2\);
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => N_58162,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_51__G2\);
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => N_58161,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_24__G2\);
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => N_58160,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_1__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP1\);
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => N_58159,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_53__G2\);
RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000010000000")
port map (
combout => N_58158,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN11_WQSTSETS\);
RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M14S2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111111")
port map (
combout => N_58157,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_10__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_7__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M11S4_RETI\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_6_RETI\);
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => N_58156,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_50__G2\);
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => N_58155,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_48__G2\);
RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN15_NOTXZYFROMD_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110010100000")
port map (
combout => N_58154,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_375__G0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(11));
RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN16_NOTXZYFROMD: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => N_58153,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(1));
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => N_58152,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_30__G2\);
\RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100111110101111")
port map (
combout => N_58151,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.UN10_U_SNNOTDB_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.TOGGLESIG\);
RETGRLFPC2_0_FPI_LDOP: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => N_58150,
dataa => \GRLFPC2_0.RIN.MK.LDOP_7\,
datab => \GRLFPC2_0.RIN.MK.LDOP_8\,
datac => \GRLFPC2_0.RIN.MK.LDOP_9\,
datad => \GRLFPC2_0.FPI.LDOP_0_X\);
RETGRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN3_NOTXZYFROMD: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000111110001111")
port map (
combout => N_58149,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_DIVMULTV\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD_A_RETI\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_173_RNIT8MM: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63),
dataa => \GRLFPC2_0.FPI.LDOP_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(63),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(63));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_EXTEND_TEMP_1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.EXTEND.TEMP_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5416\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN26_XZYBUSLSBS\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_170_RNIN8MM: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62),
dataa => \GRLFPC2_0.FPI.LDOP_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(62));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_167_RNI31MM: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
dataa => \GRLFPC2_0.FPI.LDOP_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(61));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_164_RNIT0MM: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
dataa => \GRLFPC2_0.FPI.LDOP_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(64),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(64));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_161_RNIN0MM: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
dataa => \GRLFPC2_0.FPI.LDOP_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(77));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_158_RNI3PLM: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69),
dataa => \GRLFPC2_0.FPI.LDOP_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(69),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(69));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_155_RNITOLM: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
dataa => \GRLFPC2_0.FPI.LDOP_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(68),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(68));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_152_RNINOLM: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67),
dataa => \GRLFPC2_0.FPI.LDOP_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(67),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(67));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_149_RNIQKLM: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
dataa => \GRLFPC2_0.FPI.LDOP_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(76),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(76));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_146_RNITGLM: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75),
dataa => \GRLFPC2_0.FPI.LDOP_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(75),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(75));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_143_RNINGLM: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
dataa => \GRLFPC2_0.FPI.LDOP_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(74),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(74));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_140_RNIHGLM: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73),
dataa => \GRLFPC2_0.FPI.LDOP_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(73),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(73));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_137_RNIT8LM: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
dataa => \GRLFPC2_0.FPI.LDOP_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(72),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(72));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_134_RNIN8LM: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
dataa => \GRLFPC2_0.FPI.LDOP_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(71),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(71));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIJKQ7_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_48__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_48__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0_RETI\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_RETI\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_RETI\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_RNO_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_49__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNI5KO7_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_50__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(50));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_50__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_49__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0_RETI\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_RETI\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_RETI\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_129_RNIM4LM: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70),
dataa => \GRLFPC2_0.FPI.LDOP_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(70),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(70));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M14_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M14_RETI\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M14S2_RETI\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12_RETI\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13_RETI\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_COUNTSUCCESSIVEZERO36: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_7_RETI\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_6_RETI\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_8_RETI\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_A_RETI\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_10_RNI4SOM: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100011001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_M_RETO\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_RETO\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_RNO_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_21__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(21),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_21__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_122_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122_RETI\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNI7KP7_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_24__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(24),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIBCP7_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_53__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_53__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_24__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN8_TEMP_2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000011011101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN8_TEMP_2_RETI\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(24),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN8_TEMP_2_A_RETI\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNI7SO7_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_51__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNI94P7_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_52__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_52__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_51__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0_RETI\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_RETI\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_RETI\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS_RETI\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS_2_RETI\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_115__G0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_215_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(215),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(215),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD16\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_RETI\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(215),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN25_NOTXZYFROMD_RETI\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_RETI\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD_RETI\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_216_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(216),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(216),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD15\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_RETI\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(216),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN25_NOTXZYFROMD_RETI\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_RETI\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD_RETI\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_217_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(217),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(217),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD14\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_RETI\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(217),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN25_NOTXZYFROMD_RETI\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_RETI\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD_RETI\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_218_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(218),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(218),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD13\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_13_M1_E: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_13_M1_E_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1_RETI\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN25_NOTXZYFROMD_RETI\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_13_M1_E_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD_RETI\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_13_M1_E_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010001010100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_13_M1_E_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(218),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_219_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(219),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(219),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD12\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_RETI\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(219),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN25_NOTXZYFROMD_RETI\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_RETI\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD_RETI\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_220_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(220),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(220),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD11\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_RETI\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(220),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN25_NOTXZYFROMD_RETI\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_RETI\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD_RETI\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_221_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(221),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(221),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD10\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_RETI\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(221),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN25_NOTXZYFROMD_RETI\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_RETI\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD_RETI\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_222_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(222),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(222),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD9\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_RETI\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(222),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN25_NOTXZYFROMD_RETI\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_RETI\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD_RETI\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_223_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(223),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(223),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_RETI\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(223),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN25_NOTXZYFROMD_RETI\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_RETI\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD_RETI\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_228_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(228),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(228),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_3_M1_E_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_3_M1_E_1_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(228),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN25_NOTXZYFROMD_RETI\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD_RETI\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_REP1EN_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1I\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_16__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100011001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS_2_RETI\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.UN53_SCTRL_NEW\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1I\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_0_0_3__G0_I\);
GRLFPC2_0_R_MK_BUSY_RET_RNIKO6A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.R.MK.BUSY_RET\,
dataa => RST_RETO,
datab => \GRLFPC2_0.R.MK.RST_RET_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_64_RNI45LB: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_60_RNIB2RQ: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_RETO\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_RETO\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN14_CONDITIONAL_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_58_RNI95LB: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_X_RETO\(0),
dataa => CPI_D_INST_RETO(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_55_RNIBAAN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010101000111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_0_RETO\,
dataa => CPI_D_INST_RETO(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_7_1_RETO\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_51_RNI3AAN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010101000111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_84__G0_0_RETO\,
dataa => CPI_D_INST_RETO(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_0_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47_RNIDAAN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000101011001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_78__G0_0_RETO\,
dataa => CPI_D_INST_RETO(12),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_42_RNID2RQ: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101011000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO\,
dataa => CPI_D_INST_RETO(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_2_0_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_40_RNI6AAN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000101011001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_6__G0_0_RETO\,
dataa => CPI_D_INST_RETO(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2_RETO\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_35_RNI7AAN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010101000111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_0__G0_0_RETO\,
dataa => CPI_D_INST_RETO(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_RETO\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M5_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011001000110010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5_RETI\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_12__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_11__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_13__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M2_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011001000110010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M2_RETI\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_16__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_15__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_17__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M8_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111000001110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M8_RETI\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_8__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_9__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_7__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M11_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011001000110010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M11_RETI\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_4__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_3__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_5__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M13_0_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13_0_RETI\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_8__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_9__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_7__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M12_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12_RETI\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_15__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_16__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_17__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5S4_RETI\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M12_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111111101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12_RETI\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_17__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M2S2_RETI\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5S4_1_RETI\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5S4_RETI\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M13_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011111100111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13_RETI\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_9__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M11S4_1_RETI\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M11S4_RETI\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M8S2_RETI\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M14S2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M14S2_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_10__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_7__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M11S4_RETI\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_6_RETI\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_COUNTSUCCESSIVEZERO36_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_A_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_3__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_14__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_A_S_RETI\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_COUNTSUCCESSIVEZERO36_8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_8_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_4__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_5__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_6__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_7__G2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_COUNTSUCCESSIVEZERO36_7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_7_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_2__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_10__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_15__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_17__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M5_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110011011100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5_RETI\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_12__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_11__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_13__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M8_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111010011110100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M8_RETI\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_8__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_9__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_7__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110011011100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M2_RETI\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_16__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_15__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_17__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M11_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110011011100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M11_RETI\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_4__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_3__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_5__G2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_6_M3_E: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_6_M3_E_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1_RETI\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN25_NOTXZYFROMD_RETI\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_6_M3_E_0_RETI\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD_RETI\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_95_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000111001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM_A_RETI\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_RETI\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_2_M1_E_1_RETI\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1_RETI\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_91_RNIB70Q: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001100100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_372__G1_RETO\,
datab => \GRLFPC2_0.FPI.LDOP_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(113));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_85_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_84_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_224_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(224),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(224),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD7\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_7_M3_E_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_7_M3_E_1_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(224),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1_RETI\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_225_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(225),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(225),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD6\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_6_M3_E_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010001010100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_6_M3_E_0_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(225),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_81_RNI870Q: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111111101010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
dataa => \GRLFPC2_0.FPI.LDOP_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_319__G1_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(60));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_80_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_112__G2\,
dataa => N_670,
datab => \GRLFPC2_0.FPI.LDOP_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(112));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_80_RNICLM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_112__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_78_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_111__G2\,
dataa => N_671,
datab => \GRLFPC2_0.FPI.LDOP_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(111));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_78_RNIJLM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_111__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_76_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_110__G2\,
dataa => N_672,
datab => \GRLFPC2_0.FPI.LDOP_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(110));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_76_RNIHLM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_110__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_74_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_109__G2\,
dataa => N_673,
datab => \GRLFPC2_0.FPI.LDOP_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(109));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_74_RNIFLM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_109__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_72_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_108__G2\,
dataa => N_674,
datab => \GRLFPC2_0.FPI.LDOP_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(108));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_72_RNIDLM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_108__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_70_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_107__G2\,
dataa => N_675,
datab => \GRLFPC2_0.FPI.LDOP_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(107));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_70_RNIBLM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_107__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_68_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_106__G2\,
dataa => N_676,
datab => \GRLFPC2_0.FPI.LDOP_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(106));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_68_RNIILM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_106__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_66_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_105__G2\,
dataa => N_677,
datab => \GRLFPC2_0.FPI.LDOP_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(105));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_66_RNIGLM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_105__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_64_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_104__G2\,
dataa => N_678,
datab => \GRLFPC2_0.FPI.LDOP_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(104));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_64_RNIELM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_104__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_62_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_103__G2\,
dataa => N_679,
datab => \GRLFPC2_0.FPI.LDOP_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(103));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_62_RNICLM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_103__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_60_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_102__G2\,
dataa => N_680,
datab => \GRLFPC2_0.FPI.LDOP_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(102));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_60_RNIALM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_102__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_58_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_101__G2\,
dataa => N_681,
datab => \GRLFPC2_0.FPI.LDOP_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(101));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_58_RNIHLM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_101__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_56_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_100__G2\,
dataa => N_682,
datab => \GRLFPC2_0.FPI.LDOP_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(100));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_56_RNIFLM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_100__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_54_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_99__G2\,
dataa => N_683,
datab => \GRLFPC2_0.FPI.LDOP_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(99));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_54_RNIDLM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_99__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_52_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_98__G2\,
dataa => N_684,
datab => \GRLFPC2_0.FPI.LDOP_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(98));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_52_RNIBLM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_98__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_50_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_97__G2\,
dataa => N_685,
datab => \GRLFPC2_0.FPI.LDOP_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(97));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_50_RNI9LM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_97__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_48_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_96__G2\,
dataa => N_686,
datab => \GRLFPC2_0.FPI.LDOP_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(96));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_48_RNIGLM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_96__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_46_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_95__G2\,
dataa => N_687,
datab => \GRLFPC2_0.FPI.LDOP_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(95));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_46_RNIELM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_95__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_44_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_94__G2\,
dataa => N_688,
datab => \GRLFPC2_0.FPI.LDOP_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(94));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_44_RNICLM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_94__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_43_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_93__G2\,
dataa => N_689,
datab => \GRLFPC2_0.FPI.LDOP_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(93));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_43_RNIBLM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_93__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_42_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_92__G2\,
dataa => N_690,
datab => \GRLFPC2_0.FPI.LDOP_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(92));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_42_RNIALM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_92__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_41_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_91__G2\,
dataa => N_691,
datab => \GRLFPC2_0.FPI.LDOP_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(91));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_41_RNI9LM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_91__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_40_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_90__G2\,
dataa => N_692,
datab => \GRLFPC2_0.FPI.LDOP_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(90));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_40_RNI8LM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_90__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_39_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_89__G2\,
dataa => N_693,
datab => \GRLFPC2_0.FPI.LDOP_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(89));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_39_RNIGLM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_89__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_38_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_88__G2\,
dataa => N_694,
datab => \GRLFPC2_0.FPI.LDOP_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(88));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_38_RNIFLM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_88__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_37_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_87__G2\,
dataa => N_695,
datab => \GRLFPC2_0.FPI.LDOP_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(87));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_37_RNIELM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_87__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_35_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_86__G2\,
dataa => N_696,
datab => \GRLFPC2_0.FPI.LDOP_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(86));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_35_RNICLM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_86__G2_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_33_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100110010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1_RETI\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN25_NOTXZYFROMD_RETI\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1_RETI\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD_RETI\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_4_M3_E: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_4_M3_E_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1_RETI\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN25_NOTXZYFROMD_RETI\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_4_M3_E_0_RETI\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD_RETI\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_31_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1_RETI\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN25_NOTXZYFROMD_RETI\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1_RETI\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD_RETI\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M11S4_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M11S4_1_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_4__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_3__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_5__G2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M5S4_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5S4_1_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_11__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_12__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_13__G2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M8S2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M8S2_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_8__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_7__G2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M2S2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M2S2_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_16__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_15__G2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M5S4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5S4_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_14__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_11__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_12__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_13__G2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_COUNTSUCCESSIVEZERO36_6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_6_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_9__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_8__G2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_COUNTSUCCESSIVEZERO36_A_S: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_A_S_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_16__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_13__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_12__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_11__G2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M11S4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M11S4_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_4__G2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_3__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_5__G2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_6__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_EXTEND_TEMP_1_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000111100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.EXTEND.TEMP_1_RETI\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.EXTEND.TEMP_1_A_RETI\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_58__G0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIDKP7_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_54__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNI9SP7_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_25__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(25));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_25__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_54__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN8_TEMP_2_A_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011001010111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN8_TEMP_2_A_RETI\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_227_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(227),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(227),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_4_M3_E_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010001010100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_4_M3_E_0_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(227),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_226_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(226),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(226),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_5_M3_E_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_5_M3_E_1_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(226),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1_RETI\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_229_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(229),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(229),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_2_M1_E_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_2_M1_E_1_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(229),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN25_NOTXZYFROMD_RETI\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD_RETI\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIFSP7_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_55__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_230_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(230),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(230),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_55__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_EXTEND_TEMP_1_A_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001101011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.EXTEND.TEMP_1_A_RETI\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(230),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN25_NOTXZYFROMD_RETI\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD_RETI\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_231_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(231),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(231),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN26_XZYBUSLSBS: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN26_XZYBUSLSBS_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(231),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN25_NOTXZYFROMD_RETI\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_8__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_SUB_REP2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000110110001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP2_RETI\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_58__G0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN16_NOTXZYFROMD: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN15_NOTXZYFROMD_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110010100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_375__G0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN15_NOTXZYFROMD: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011110010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1_RETI\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_95_RNO_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100110010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1_RETI\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN25_NOTXZYFROMD_RETI\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1_RETI\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD_RETI\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_59__G0_XX_MM\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_59__G0_YY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_59__G0_XX\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_29_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101000100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G_32\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_23_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001110100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G_32\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_20_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_6\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_C\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_26_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_C\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_17_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_C\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_14_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_C\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNITJO7_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_10__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_COUNTSUCCESSIVEZERO36_7_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_2__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIBCQ7_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_17__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNI7SP7_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_15__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIBPDF_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_8__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIDPDF_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_9__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNI5KP7_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_14__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(14));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNI3CP7_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_13__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNI14P7_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_12__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNI94Q7_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_16__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNIVRO7_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_11__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNI9PDF_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_7__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNI3PDF_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_4__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNI5PDF_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_5__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNI7PDF_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_6__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNI1PDF_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_3__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_114_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_114__G0\,
dataa => \GRLFPC2_0.FPI.LDOP_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_3\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(114));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN38_SHDVAR_3_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_57__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(57));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_1_RNILJ4A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2_REP1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN25_NOTXZYFROMD\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_33_RNIS0E21: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_80__G0_A_RETO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_RETO\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_C_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_LI_19_M_RETO\(79));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_30_RNI363E1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_1_RETO\,
dataa => CPI_D_INST_RETO(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_I_M_RETO\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_26_RNIB63E1_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_1_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_6__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_23_RNI463E1_7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_4_0_RETO\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_20_RNI70DC1_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_U_RETO\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_6_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_84__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_17_RNII63E1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_2_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_78__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_14_RNI663E1_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_7_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_0__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_12_RNIPRP02: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_M_RETO\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_8_RNIR9B12_5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_RETO\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_C_RETO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D_RETO\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_83__G0_1_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_4_RNIN52O1_4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.FPINST_I_M_X_RETO\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_80__G0_A_RETO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN3_NOTXZYFROMD: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000111110001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_DIVMULTV\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD_A_RETI\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(12),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN25_NOTXZYFROMD: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN25_NOTXZYFROMD_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_374__G0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(12),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN16_NOTXZYFROMD_REP1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_9__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN15_NOTXZYFROMD_0_REP1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110010100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_375__G0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_RNITODF_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_1__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_REP0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(14),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_14__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHEN_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_1__G2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_16__G2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN3_NOTXZYFROMD_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001101011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD_A_RETI\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(14),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(1));
\GRLFPC2_0_R_FSR_CEXC_RNO_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.R.FSR.CEXC_1_0_4__G1\,
dataa => \GRLFPC2_0.COMB.V.FSR.CEXC_1_2\(4),
datab => \GRLFPC2_0.COMB.V.FSR.CEXC_1_1_X\(4),
datac => \GRLFPC2_0.COMB.V.FSR.CEXC_1_SN_M3\);
\GRLFPC2_0_R_FSR_CEXC_RNO_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.R.FSR.CEXC_1_0_3__G1\,
dataa => \GRLFPC2_0.COMB.V.FSR.CEXC_1_2\(3),
datab => \GRLFPC2_0.COMB.V.FSR.CEXC_1_1_X\(3),
datac => \GRLFPC2_0.COMB.V.FSR.CEXC_1_SN_M3\);
\GRLFPC2_0_R_FSR_CEXC_RNO_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.R.FSR.CEXC_1_0_2__G1\,
dataa => \GRLFPC2_0.COMB.V.FSR.CEXC_1_2\(2),
datab => \GRLFPC2_0.COMB.V.FSR.CEXC_1_1_X\(2),
datac => \GRLFPC2_0.COMB.V.FSR.CEXC_1_SN_M3\);
\GRLFPC2_0_R_FSR_CEXC_RNO_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.R.FSR.CEXC_1_0_1__G1\,
dataa => \GRLFPC2_0.COMB.V.FSR.CEXC_1_2\(1),
datab => \GRLFPC2_0.COMB.V.FSR.CEXC_1_1_X\(1),
datac => \GRLFPC2_0.COMB.V.FSR.CEXC_1_SN_M3\);
\GRLFPC2_0_R_FSR_CEXC_RNO_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.R.FSR.CEXC_1_0_0__G1\,
dataa => \GRLFPC2_0.COMB.V.FSR.CEXC_1_2\(0),
datab => \GRLFPC2_0.COMB.V.FSR.CEXC_1_1_X\(0),
datac => \GRLFPC2_0.COMB.V.FSR.CEXC_1_SN_M3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_257_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(257),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\(257),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\(257),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_256_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(256),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\(256),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\(256),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_255_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(255),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\(255),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\(255),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_254_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(254),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\(254),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\(254),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_253_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(253),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\(253),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\(253),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_252_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(252),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\(252),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\(252),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_251_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(251),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\(251),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\(251),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_250_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(250),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\(250),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\(250),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_244_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__G0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_33\(244),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__G1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_243_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_243__G0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_33\(243),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_243__G1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_242_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_242__G0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_33\(242),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_242__G1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_241_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_241__G0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_33\(241),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_241__G1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_240_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_240__G0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_33\(240),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_240__G1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_239_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_239__G0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_33\(239),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_239__G1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_238_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_238__G0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_33\(238),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_238__G1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_237_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_237__G0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_33\(237),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_237__G1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_172_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(172),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_14\(172));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_171_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(171),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_14\(171));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_142_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(142),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD31\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_14\(142));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_141_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(141),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD32\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_14\(141));
\GRLFPC2_0_R_I_RES_RNO_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.COMB.V.I.RES_1\(63),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.SIGNRESULT\,
datab => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2\,
datac => \GRLFPC2_0.COMB.V.I.RES_6_X\(63));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2S2_REP3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.WQSCTRL_0_3947\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2S2_REP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.WQSCTRL_0_3947\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2S2_REP1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.WQSCTRL_0_3947\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_SUB_REP1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110110001101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_REP2_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_A\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_REP1_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_A\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_REP3_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110110001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19_3_0_.M4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_SN_M3_E\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_REP2_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110110001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19_3_0_.M4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_SN_M3_E\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_REP1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110110001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19_3_0_.M4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_SN_M3_E\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_REP2_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_SN_M3_E\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19_3_0_.M3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_REP1_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_SN_M3_E\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19_3_0_.M3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA_REP1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_0\,
datac => \GRLFPC2_0.FPI.LDOP_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SS0_REP1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111000010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLBREGXZ.UN4_XZBREGLOADEN\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.WQSCTRL_0\(67),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_REP2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_SN_M3_E\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19_3_0_.M2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_REP1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_SN_M3_E\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19_3_0_.M2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001100000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_UN10_SELECTEDMIPTR: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CONDMUXMULXFF.UN4_NOTSQRTLFTCC\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_D: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001111110001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CONDMUXMULXFF.UN4_NOTSQRTLFTCC\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14_141_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110000001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_14\(141),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(143),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_T_3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14_172_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_14\(172),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.SELECTQUOBITS.NOTDIVC\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD57\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011001111001001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(10),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_7_A\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A28_0_S_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111011110100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_0_S\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_0_S\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80));
\GRLFPC2_0_FPI_OP2_X_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(40),
dataa => N_710,
datab => N_646,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(39),
dataa => N_709,
datab => N_645,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(51),
dataa => N_721,
datab => N_657,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(50),
dataa => N_720,
datab => N_656,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(48),
dataa => N_718,
datab => N_654,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(45),
dataa => N_715,
datab => N_651,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(58),
dataa => N_728,
datab => N_664,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(55),
dataa => N_725,
datab => N_661,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(52),
dataa => N_722,
datab => N_658,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(36),
dataa => N_706,
datab => N_642,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(33),
dataa => N_703,
datab => N_639,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(32),
dataa => N_702,
datab => N_638,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(34),
dataa => N_704,
datab => N_640,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(35),
dataa => N_705,
datab => N_641,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(37),
dataa => N_707,
datab => N_643,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(59),
dataa => N_729,
datab => N_665,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(60),
dataa => N_730,
datab => N_666,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(61),
dataa => N_731,
datab => N_667,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(62),
dataa => N_732,
datab => N_668,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(53),
dataa => N_723,
datab => N_659,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(54),
dataa => N_724,
datab => N_660,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(56),
dataa => N_726,
datab => N_662,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(57),
dataa => N_727,
datab => N_663,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(46),
dataa => N_716,
datab => N_652,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(47),
dataa => N_717,
datab => N_653,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(49),
dataa => N_719,
datab => N_655,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(38),
dataa => N_708,
datab => N_644,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(41),
dataa => N_711,
datab => N_647,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(42),
dataa => N_712,
datab => N_648,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(43),
dataa => N_713,
datab => N_649,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP2_X_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(44),
dataa => N_714,
datab => N_650,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
GRLFPC2_0_COMB_FPDECODE_FPOP3_0_A2_1_X_RNIL1DI: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110111011101")
port map (
combout => \GRLFPC2_0.COMB.RS1_1_SN_M2_I_X\,
dataa => N_17,
datab => \GRLFPC2_0.COMB.RS1_1_SN_M2_I_A2\);
\GRLFPC2_0_COMB_RS1_1_0_X_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.RS1_1_0_X\(3),
dataa => N_17,
datab => N_74,
datac => \GRLFPC2_0.R.A.RS1\(3));
GRLFPC2_0_COMB_FPDECODE_FPOP3_0_A2_1_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.COMB.FPDECODE.FPOP3_0_A2_1_X\,
dataa => N_77,
datab => N_80);
GRLFPC2_0_RS1V_0_SQMUXA_1_0_A2_3_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.RS1V_0_SQMUXA_1_0_A2_3_X\,
dataa => N_70,
datab => N_69);
\GRLFPC2_0_COMB_DBGDATA_4_0_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(1),
dataa => N_405,
datab => N_671,
datac => N_607);
\GRLFPC2_0_COMB_DBGDATA_4_0_X_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(16),
dataa => N_405,
datab => N_686,
datac => N_622);
\GRLFPC2_0_FPI_OP1_X_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(45),
dataa => N_683,
datab => N_619,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_FPI_OP1_X_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(48),
dataa => N_686,
datab => N_622,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_COMB_DBGDATA_4_0_X_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(13),
dataa => N_405,
datab => N_683,
datac => N_619);
GRLFPC2_0_R_MK_BUSY_RET_2_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.R.MK.BUSY_RET_2_0_0_A2_0_G0_X\,
dataa => N_8,
datab => \GRLFPC2_0.R.MK.BUSY_RET_5\);
GRLFPC2_0_R_X_FPOP_RNINRLL: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
dataa => N_17,
datab => \GRLFPC2_0.R.I.RDD_0_0_G1_0_8238_I_O4\);
GRLFPC2_0_COMB_WREN12_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.COMB.WREN12_X\,
dataa => N_366,
datab => N_365);
GRLFPC2_0_COMB_UN3_HOLDN_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC2_0.COMB.UN3_HOLDN_X\,
dataa => N_160,
datab => N_161);
GRLFPC2_0_COMB_UN1_FPCI_2_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC2_0.COMB.UN1_FPCI_2_X\,
dataa => N_229,
datab => N_230);
GRLFPC2_0_COMB_UN1_FPCI_1_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC2_0.COMB.UN1_FPCI_1_X\,
dataa => N_298,
datab => N_299);
GRLFPC2_0_R_MK_HOLDN1_0_I_A2_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.R.MK.HOLDN1_0_I_A2_X\,
dataa => N_8,
datab => \GRLFPC2_0.R.MK.RST2\);
GRLFPC2_0_R_MK_HOLDN2_RNIRLU6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.R.MK.BUSY_RET_3_0_0_A2_X\,
dataa => N_8,
datab => \GRLFPC2_0.R.MK.HOLDN2\);
\GRLFPC2_0_COMB_RS1_1_0_X_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.RS1_1_0_X\(4),
dataa => N_17,
datab => N_75,
datac => \GRLFPC2_0.R.A.RS1\(4));
GRLFPC2_0_R_I_PC_RET_60_RNI7KV4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
dataa => N_17,
datab => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_FPI_OP1_X_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(59),
dataa => N_697,
datab => N_633,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_COMB_WRDATA_4_X_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(26),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(26),
datac => \GRLFPC2_0.R.I.RES\(55));
\GRLFPC2_0_COMB_WRDATA_4_X_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(41),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(41),
datac => \GRLFPC2_0.R.I.RES\(38));
\GRLFPC2_0_COMB_WRDATA_4_X_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(58),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(58),
datac => \GRLFPC2_0.R.I.RES\(55));
\GRLFPC2_0_COMB_DBGDATA_4_0_X_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(11),
dataa => N_405,
datab => N_681,
datac => N_617);
\GRLFPC2_0_COMB_DBGDATA_4_0_X_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(24),
dataa => N_405,
datab => N_694,
datac => N_630);
\GRLFPC2_0_COMB_DBGDATA_4_0_X_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(27),
dataa => N_405,
datab => N_697,
datac => N_633);
\GRLFPC2_0_COMB_V_FSR_FCC_1_1_X_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.FCC_1_1_X\(0),
dataa => N_380,
datab => CPO_CCZ(0),
datac => \GRLFPC2_0.V.FSR.NONSTD_0_SQMUXA_6_X\);
\GRLFPC2_0_COMB_V_FSR_FCC_1_1_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.FCC_1_1_X\(1),
dataa => N_381,
datab => CPO_CCZ(1),
datac => \GRLFPC2_0.V.FSR.NONSTD_0_SQMUXA_6_X\);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_1_X_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_1_X\(0),
dataa => N_370,
datab => \GRLFPC2_0.R.FSR.CEXC\(0),
datac => \GRLFPC2_0.V.FSR.CEXC_3_SQMUXA\);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_1_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_1_X\(2),
dataa => N_372,
datab => \GRLFPC2_0.R.FSR.CEXC\(2),
datac => \GRLFPC2_0.V.FSR.CEXC_3_SQMUXA\);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_1_X_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_1_X\(4),
dataa => N_374,
datab => \GRLFPC2_0.R.FSR.CEXC\(4),
datac => \GRLFPC2_0.V.FSR.CEXC_3_SQMUXA\);
\GRLFPC2_0_FPI_OP1_X_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(32),
dataa => N_670,
datab => N_606,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_FPI_OP1_X_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(36),
dataa => N_674,
datab => N_610,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_FPI_OP1_X_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(37),
dataa => N_675,
datab => N_611,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_FPI_OP1_X_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(40),
dataa => N_678,
datab => N_614,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_FPI_OP1_X_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(42),
dataa => N_680,
datab => N_616,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_FPI_OP1_X_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(43),
dataa => N_681,
datab => N_617,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_FPI_OP1_X_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(50),
dataa => N_688,
datab => N_624,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_FPI_OP1_X_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(55),
dataa => N_693,
datab => N_629,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_FPI_OP1_X_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(56),
dataa => N_694,
datab => N_630,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_FPI_OP1_X_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(57),
dataa => N_695,
datab => N_631,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_FPI_OP1_X_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(62),
dataa => N_700,
datab => N_636,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_FPI_OP1_X_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(63),
dataa => N_701,
datab => N_637,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_COMB_RS1_1_0_X_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.RS1_1_0_X\(0),
dataa => N_17,
datab => N_71,
datac => \GRLFPC2_0.R.A.RS1\(0));
\GRLFPC2_0_COMB_RS1_1_0_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.RS1_1_0_X\(1),
dataa => N_17,
datab => N_72,
datac => \GRLFPC2_0.R.A.RS1\(1));
\GRLFPC2_0_COMB_RS1_1_0_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.RS1_1_0_X\(2),
dataa => N_17,
datab => N_73,
datac => \GRLFPC2_0.R.A.RS1\(2));
\GRLFPC2_0_FPI_OP2_X_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP2_X\(63),
dataa => N_733,
datab => N_669,
datac => \GRLFPC2_0.COMB.UN1_FPCI_4\);
\GRLFPC2_0_FPI_OP1_X_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(46),
dataa => N_684,
datab => N_620,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_COMB_WRADDR_5_X_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.WRADDR_5_X\(0),
dataa => \GRLFPC2_0.WRADDR_1_SQMUXA\,
datab => N_358,
datac => \GRLFPC2_0.R.I.INST\(25));
\GRLFPC2_0_COMB_DBGDATA_4_0_X_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(14),
dataa => N_405,
datab => N_684,
datac => N_620);
\GRLFPC2_0_FPI_OP1_X_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(39),
dataa => N_677,
datab => N_613,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_COMB_DBGDATA_4_0_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(2),
dataa => N_405,
datab => N_672,
datac => N_608);
\GRLFPC2_0_COMB_DBGDATA_4_0_X_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(7),
dataa => N_405,
datab => N_677,
datac => N_613);
\GRLFPC2_0_COMB_DBGDATA_4_0_X_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(9),
dataa => N_405,
datab => N_679,
datac => N_615);
\GRLFPC2_0_FPI_OP1_X_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(33),
dataa => N_671,
datab => N_607,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_FPI_OP1_X_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(34),
dataa => N_672,
datab => N_608,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_FPI_OP1_X_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(35),
dataa => N_673,
datab => N_609,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_FPI_OP1_X_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(41),
dataa => N_679,
datab => N_615,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_FPI_OP1_X_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(44),
dataa => N_682,
datab => N_618,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_FPI_OP1_X_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(47),
dataa => N_685,
datab => N_621,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_FPI_OP1_X_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(49),
dataa => N_687,
datab => N_623,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_FPI_OP1_X_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(51),
dataa => N_689,
datab => N_625,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_FPI_OP1_X_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(52),
dataa => N_690,
datab => N_626,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_FPI_OP1_X_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(53),
dataa => N_691,
datab => N_627,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_FPI_OP1_X_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(54),
dataa => N_692,
datab => N_628,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_FPI_OP1_X_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(60),
dataa => N_698,
datab => N_634,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_FPI_OP1_X_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(61),
dataa => N_699,
datab => N_635,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_COMB_WRADDR_5_I_M2_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.WRADDR_5_I_M2_X\(1),
dataa => \GRLFPC2_0.WRADDR_1_SQMUXA\,
datab => N_359,
datac => \GRLFPC2_0.R.I.INST\(26));
\GRLFPC2_0_COMB_WRADDR_5_I_M2_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.WRADDR_5_I_M2_X\(2),
dataa => \GRLFPC2_0.WRADDR_1_SQMUXA\,
datab => N_360,
datac => \GRLFPC2_0.R.I.INST\(27));
\GRLFPC2_0_COMB_WRADDR_5_I_M2_X_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.WRADDR_5_I_M2_X\(3),
dataa => \GRLFPC2_0.WRADDR_1_SQMUXA\,
datab => N_361,
datac => \GRLFPC2_0.R.I.INST\(28));
\GRLFPC2_0_COMB_WRDATA_4_X_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(54),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(54),
datac => \GRLFPC2_0.R.I.RES\(51));
\GRLFPC2_0_COMB_DBGDATA_4_0_X_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(3),
dataa => N_405,
datab => N_673,
datac => N_609);
\GRLFPC2_0_COMB_DBGDATA_4_0_X_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(22),
dataa => N_405,
datab => N_692,
datac => N_628);
\GRLFPC2_0_COMB_WRDATA_4_X_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(4),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(4),
datac => \GRLFPC2_0.R.I.RES\(33));
\GRLFPC2_0_COMB_WRDATA_4_X_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(29),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(29),
datac => \GRLFPC2_0.R.I.RES\(58));
\GRLFPC2_0_COMB_WRDATA_4_X_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(36),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(36),
datac => \GRLFPC2_0.R.I.RES\(33));
\GRLFPC2_0_COMB_WRDATA_4_X_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(61),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(61),
datac => \GRLFPC2_0.R.I.RES\(58));
\GRLFPC2_0_COMB_WRDATA_4_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(1),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(1),
datac => \GRLFPC2_0.R.I.RES\(30));
\GRLFPC2_0_COMB_WRDATA_4_X_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(22),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(22),
datac => \GRLFPC2_0.R.I.RES\(51));
\GRLFPC2_0_COMB_WRDATA_4_X_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(33),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(33),
datac => \GRLFPC2_0.R.I.RES\(30));
\GRLFPC2_0_COMB_V_FSR_CEXC_1_1_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_1_X\(1),
dataa => N_371,
datab => \GRLFPC2_0.R.FSR.CEXC\(1),
datac => \GRLFPC2_0.V.FSR.CEXC_3_SQMUXA\);
\GRLFPC2_0_COMB_WRDATA_4_X_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(15),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(15),
datac => \GRLFPC2_0.R.I.RES\(44));
\GRLFPC2_0_COMB_WRDATA_4_X_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(18),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(18),
datac => \GRLFPC2_0.R.I.RES\(47));
\GRLFPC2_0_COMB_WRDATA_4_X_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(21),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(21),
datac => \GRLFPC2_0.R.I.RES\(50));
\GRLFPC2_0_COMB_WRDATA_4_X_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(47),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(47),
datac => \GRLFPC2_0.R.I.RES\(44));
\GRLFPC2_0_COMB_WRDATA_4_X_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(50),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(50),
datac => \GRLFPC2_0.R.I.RES\(47));
\GRLFPC2_0_COMB_WRDATA_4_X_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(53),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(53),
datac => \GRLFPC2_0.R.I.RES\(50));
\GRLFPC2_0_COMB_WRDATA_4_X_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(12),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(12),
datac => \GRLFPC2_0.R.I.RES\(41));
\GRLFPC2_0_COMB_WRDATA_4_X_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(24),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(24),
datac => \GRLFPC2_0.R.I.RES\(53));
\GRLFPC2_0_COMB_WRDATA_4_X_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(32),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(32),
datac => \GRLFPC2_0.R.I.RES\(29));
\GRLFPC2_0_COMB_WRDATA_4_X_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(44),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(44),
datac => \GRLFPC2_0.R.I.RES\(41));
\GRLFPC2_0_COMB_WRDATA_4_X_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(56),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(56),
datac => \GRLFPC2_0.R.I.RES\(53));
\GRLFPC2_0_COMB_WRADDR_5_X_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.WRADDR_5_X\(4),
dataa => \GRLFPC2_0.WRADDR_1_SQMUXA\,
datab => N_362,
datac => \GRLFPC2_0.R.I.INST\(29));
\GRLFPC2_0_COMB_DBGDATA_4_0_X_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(23),
dataa => N_405,
datab => N_693,
datac => N_629);
\GRLFPC2_0_FPI_OP1_X_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(38),
dataa => N_676,
datab => N_612,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_COMB_WRDATA_4_X_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(5),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(5),
datac => \GRLFPC2_0.R.I.RES\(34));
\GRLFPC2_0_COMB_WRDATA_4_X_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(6),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(6),
datac => \GRLFPC2_0.R.I.RES\(35));
\GRLFPC2_0_COMB_WRDATA_4_X_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(37),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(37),
datac => \GRLFPC2_0.R.I.RES\(34));
\GRLFPC2_0_COMB_WRDATA_4_X_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(38),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(38),
datac => \GRLFPC2_0.R.I.RES\(35));
\GRLFPC2_0_COMB_DBGDATA_4_0_X_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(5),
dataa => N_405,
datab => N_675,
datac => N_611);
\GRLFPC2_0_COMB_DBGDATA_4_0_X_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(6),
dataa => N_405,
datab => N_676,
datac => N_612);
\GRLFPC2_0_COMB_DBGDATA_4_0_X_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(8),
dataa => N_405,
datab => N_678,
datac => N_614);
\GRLFPC2_0_FPI_OP1_X_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.FPI.OP1_X\(58),
dataa => N_696,
datab => N_632,
datac => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_COMB_WRDATA_4_X_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(25),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(25),
datac => \GRLFPC2_0.R.I.RES\(54));
\GRLFPC2_0_COMB_WRDATA_4_X_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(27),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(27),
datac => \GRLFPC2_0.R.I.RES\(56));
\GRLFPC2_0_COMB_WRDATA_4_X_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(30),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(30),
datac => \GRLFPC2_0.R.I.RES\(59));
\GRLFPC2_0_COMB_WRDATA_4_X_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(57),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(57),
datac => \GRLFPC2_0.R.I.RES\(54));
\GRLFPC2_0_COMB_WRDATA_4_X_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(59),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(59),
datac => \GRLFPC2_0.R.I.RES\(56));
\GRLFPC2_0_COMB_WRDATA_4_X_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(62),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(62),
datac => \GRLFPC2_0.R.I.RES\(59));
\GRLFPC2_0_COMB_V_FSR_TEM_1_0_X_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.TEM_1_0_X\(0),
dataa => N_393,
datab => \GRLFPC2_0.R.FSR.TEM\(0),
datac => \GRLFPC2_0.V.FSR.NONSTD_0_SQMUXA_6_X\);
\GRLFPC2_0_COMB_V_FSR_TEM_1_0_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.TEM_1_0_X\(2),
dataa => N_395,
datab => \GRLFPC2_0.R.FSR.TEM\(2),
datac => \GRLFPC2_0.V.FSR.NONSTD_0_SQMUXA_6_X\);
\GRLFPC2_0_COMB_V_FSR_TEM_1_0_X_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.TEM_1_0_X\(3),
dataa => N_396,
datab => \GRLFPC2_0.R.FSR.TEM\(3),
datac => \GRLFPC2_0.V.FSR.NONSTD_0_SQMUXA_6_X\);
\GRLFPC2_0_COMB_V_FSR_TEM_1_0_X_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.TEM_1_0_X\(4),
dataa => N_397,
datab => \GRLFPC2_0.R.FSR.TEM\(4),
datac => \GRLFPC2_0.V.FSR.NONSTD_0_SQMUXA_6_X\);
\GRLFPC2_0_COMB_V_FSR_RD_1_0_X_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.RD_1_0_X\(0),
dataa => N_400,
datab => \GRLFPC2_0.R.FSR.RD\(0),
datac => \GRLFPC2_0.V.FSR.NONSTD_0_SQMUXA_6_X\);
\GRLFPC2_0_COMB_V_FSR_RD_1_0_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.RD_1_0_X\(1),
dataa => N_401,
datab => \GRLFPC2_0.R.FSR.RD\(1),
datac => \GRLFPC2_0.V.FSR.NONSTD_0_SQMUXA_6_X\);
\GRLFPC2_0_COMB_DBGDATA_4_0_X_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(0),
dataa => N_405,
datab => N_670,
datac => N_606);
\GRLFPC2_0_COMB_DBGDATA_4_0_X_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(4),
dataa => N_405,
datab => N_674,
datac => N_610);
\GRLFPC2_0_COMB_DBGDATA_4_0_X_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(10),
dataa => N_405,
datab => N_680,
datac => N_616);
\GRLFPC2_0_COMB_DBGDATA_4_0_X_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(25),
dataa => N_405,
datab => N_695,
datac => N_631);
\GRLFPC2_0_COMB_DBGDATA_4_0_X_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(26),
dataa => N_405,
datab => N_696,
datac => N_632);
\GRLFPC2_0_COMB_DBGDATA_4_0_X_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(30),
dataa => N_405,
datab => N_700,
datac => N_636);
\GRLFPC2_0_COMB_DBGDATA_4_0_X_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(31),
dataa => N_405,
datab => N_701,
datac => N_637);
\GRLFPC2_0_COMB_WRDATA_4_X_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(8),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(8),
datac => \GRLFPC2_0.R.I.RES\(37));
\GRLFPC2_0_COMB_WRDATA_4_X_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(11),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(11),
datac => \GRLFPC2_0.R.I.RES\(40));
\GRLFPC2_0_COMB_WRDATA_4_X_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(14),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(14),
datac => \GRLFPC2_0.R.I.RES\(43));
\GRLFPC2_0_COMB_WRDATA_4_X_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(17),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(17),
datac => \GRLFPC2_0.R.I.RES\(46));
\GRLFPC2_0_COMB_WRDATA_4_X_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(20),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(20),
datac => \GRLFPC2_0.R.I.RES\(49));
\GRLFPC2_0_COMB_WRDATA_4_X_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(23),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(23),
datac => \GRLFPC2_0.R.I.RES\(52));
\GRLFPC2_0_COMB_WRDATA_4_X_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(31),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(31),
datac => \GRLFPC2_0.R.I.RES\(63));
\GRLFPC2_0_COMB_WRDATA_4_X_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(40),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(40),
datac => \GRLFPC2_0.R.I.RES\(37));
\GRLFPC2_0_COMB_WRDATA_4_X_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(43),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(43),
datac => \GRLFPC2_0.R.I.RES\(40));
\GRLFPC2_0_COMB_WRDATA_4_X_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(46),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(46),
datac => \GRLFPC2_0.R.I.RES\(43));
\GRLFPC2_0_COMB_WRDATA_4_X_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(49),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(49),
datac => \GRLFPC2_0.R.I.RES\(46));
\GRLFPC2_0_COMB_WRDATA_4_X_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(52),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(52),
datac => \GRLFPC2_0.R.I.RES\(49));
\GRLFPC2_0_COMB_WRDATA_4_X_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(55),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(55),
datac => \GRLFPC2_0.R.I.RES\(52));
\GRLFPC2_0_WRDATA_0_X_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(63),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_401,
datac => \GRLFPC2_0.R.I.RES\(63));
\GRLFPC2_0_COMB_WRDATA_4_X_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(13),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(13),
datac => \GRLFPC2_0.R.I.RES\(42));
\GRLFPC2_0_COMB_WRDATA_4_X_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(16),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(16),
datac => \GRLFPC2_0.R.I.RES\(45));
\GRLFPC2_0_COMB_WRDATA_4_X_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(19),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(19),
datac => \GRLFPC2_0.R.I.RES\(48));
\GRLFPC2_0_COMB_WRDATA_4_X_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(28),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(28),
datac => \GRLFPC2_0.R.I.RES\(57));
\GRLFPC2_0_COMB_WRDATA_4_X_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(45),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(45),
datac => \GRLFPC2_0.R.I.RES\(42));
\GRLFPC2_0_COMB_WRDATA_4_X_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(48),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(48),
datac => \GRLFPC2_0.R.I.RES\(45));
\GRLFPC2_0_COMB_WRDATA_4_X_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(51),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(51),
datac => \GRLFPC2_0.R.I.RES\(48));
GRLFPC2_0_COMB_V_FSR_NONSTD_1_0_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.NONSTD_1_0_X\,
dataa => N_392,
datab => \GRLFPC2_0.R.FSR.NONSTD\,
datac => \GRLFPC2_0.V.FSR.NONSTD_0_SQMUXA_6_X\);
\GRLFPC2_0_COMB_WRDATA_4_X_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(7),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(7),
datac => \GRLFPC2_0.R.I.RES\(36));
\GRLFPC2_0_COMB_WRDATA_4_X_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(9),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(9),
datac => \GRLFPC2_0.R.I.RES\(38));
\GRLFPC2_0_COMB_WRDATA_4_X_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(39),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(39),
datac => \GRLFPC2_0.R.I.RES\(36));
\GRLFPC2_0_COMB_WRDATA_4_X_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(60),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(60),
datac => \GRLFPC2_0.R.I.RES\(57));
\GRLFPC2_0_COMB_WRDATA_4_X_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(0),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(0),
datac => \GRLFPC2_0.R.I.RES\(29));
\GRLFPC2_0_COMB_WRDATA_4_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(2),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(2),
datac => \GRLFPC2_0.R.I.RES\(31));
\GRLFPC2_0_COMB_WRDATA_4_X_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(3),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(3),
datac => \GRLFPC2_0.R.I.RES\(32));
\GRLFPC2_0_COMB_WRDATA_4_X_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(10),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(10),
datac => \GRLFPC2_0.R.I.RES\(39));
\GRLFPC2_0_COMB_WRDATA_4_X_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(34),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(34),
datac => \GRLFPC2_0.R.I.RES\(31));
\GRLFPC2_0_COMB_WRDATA_4_X_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(35),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(35),
datac => \GRLFPC2_0.R.I.RES\(32));
\GRLFPC2_0_COMB_WRDATA_4_X_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.COMB.WRDATA_4_X\(42),
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.R.I.RES\(42),
datac => \GRLFPC2_0.R.I.RES\(39));
\GRLFPC2_0_COMB_V_FSR_TEM_1_0_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.TEM_1_0_X\(1),
dataa => N_394,
datab => \GRLFPC2_0.R.FSR.TEM\(1),
datac => \GRLFPC2_0.V.FSR.NONSTD_0_SQMUXA_6_X\);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_1_X_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_1_X\(3),
dataa => N_373,
datab => \GRLFPC2_0.R.FSR.CEXC\(3),
datac => \GRLFPC2_0.V.FSR.CEXC_3_SQMUXA\);
GRLFPC2_0_COMB_UN31_DEBUG_UNIT_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
dataa => N_403,
datab => N_404);
\GRLFPC2_0_COMB_RS1_1_1_X_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.COMB.RS1_1_1_X\(0),
dataa => \GRLFPC2_0.RS1V_0_SQMUXA_0_A2_X\,
datab => N_82);
GRLFPC2_0_RS1V_0_SQMUXA_1_0_A2_2_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.RS1V_0_SQMUXA_1_0_A2_2_X\,
dataa => N_67,
datab => N_68);
GRLFPC2_0_RS1V_0_SQMUXA_1_0_A2_1_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.RS1V_0_SQMUXA_1_0_A2_1_X\,
dataa => N_76,
datab => N_66);
GRLFPC2_0_COMB_V_E_STDATA2_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
dataa => N_159,
datab => N_158);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW_6_0_0__G2_0_X\,
dataa => N_68,
datab => N_64);
GRLFPC2_0_R_A_LD_RNO_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC2_0.N_939_I_I_2_0_X\,
dataa => N_18,
datab => N_91);
GRLFPC2_0_COMB_LOCK_1_1_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.COMB.LOCK_1_1_X\,
dataa => N_92,
datab => \GRLFPC2_0.N_939_I_I_A2\);
GRLFPC2_0_COMB_RDD_1_M14_0_A2_2_2_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.COMB.RDD_1.M14_0_A2_2_2_X\,
dataa => N_70,
datab => N_68);
\GRLFPC2_0_COMB_DBGDATA_4_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(1),
dataa => N_404,
datab => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(1),
datac => \GRLFPC2_0.R.FSR.CEXC\(1));
\GRLFPC2_0_COMB_DBGDATA_4_X_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(16),
dataa => N_404,
datab => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(16),
datac => \GRLFPC2_0.R.FSR.FTT\(2));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(19),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(19),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(19));
GRLFPC2_0_R_A_FPOP_RNIE2QG: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC2_0.R.E.FPOP_0_0_G1_X\,
dataa => N_161,
datab => N_160,
datac => \GRLFPC2_0.R.A.FPOP\);
GRLFPC2_0_R_E_LD_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC2_0.R.E.LD_0_0_G1_X\,
dataa => N_161,
datab => N_160,
datac => \GRLFPC2_0.R.A.LD\);
GRLFPC2_0_R_M_FPOP_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC2_0.R.M.FPOP_0_0_G1_X\,
dataa => N_230,
datab => N_229,
datac => \GRLFPC2_0.R.E.FPOP\);
GRLFPC2_0_R_M_LD_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC2_0.R.M.LD_0_0_G1_X\,
dataa => N_230,
datab => N_229,
datac => \GRLFPC2_0.R.E.LD\);
GRLFPC2_0_R_X_FPOP_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC2_0.R.X.FPOP_0_0_G1_X\,
dataa => N_299,
datab => N_298,
datac => \GRLFPC2_0.R.M.FPOP\);
GRLFPC2_0_R_X_LD_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC2_0.R.X.LD_0_0_G1_X\,
dataa => N_299,
datab => N_298,
datac => \GRLFPC2_0.R.M.LD\);
GRLFPC2_0_COMB_FPDECODE_ST_0_A2_0_A2_0_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC2_0.COMB.FPDECODE.ST_0_A2_0_A2_0_X\,
dataa => N_81,
datab => N_79,
datac => N_78);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_X_81_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_X\(81),
dataa => N_701,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.FPI.OP1_X\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_X_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1_X\(23),
dataa => N_733,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.FPI.OP2_X\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_X_83_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_X\(83),
dataa => N_699,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.FPI.OP1_X\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_X_82_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_X\(82),
dataa => N_700,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.FPI.OP1_X\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_X_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1_X\(24),
dataa => N_732,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.FPI.OP2_X\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_X_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1_X\(25),
dataa => N_731,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.FPI.OP2_X\(32));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(23),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(23),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(23));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(24),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(24),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(24));
\GRLFPC2_0_COMB_DBGDATA_4_X_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(11),
dataa => N_404,
datab => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(11),
datac => CPO_CCZ(1));
\GRLFPC2_0_COMB_DBGDATA_4_X_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(24),
dataa => N_404,
datab => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(24),
datac => \GRLFPC2_0.R.FSR.TEM\(1));
\GRLFPC2_0_COMB_DBGDATA_4_X_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(27),
dataa => N_404,
datab => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(27),
datac => \GRLFPC2_0.R.FSR.TEM\(4));
\GRLFPC2_0_WRDATA_0_X_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(26),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_396,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(26));
\GRLFPC2_0_WRDATA_0_X_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(41),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_379,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(41));
\GRLFPC2_0_WRDATA_0_X_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(58),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_396,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(58));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(2),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(2),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(2));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(3),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(3),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(3));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(4),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(4),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(4));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(5),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(5),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(5));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(6),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(6),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(6));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(28),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(28),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(28));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(17),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(17),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(17));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(18),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(18),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(18));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(25),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(25),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(25));
\GRLFPC2_0_COMB_DBGDATA_4_X_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(14),
dataa => N_404,
datab => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(14),
datac => \GRLFPC2_0.R.FSR.FTT\(0));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(26),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(26),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(26));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(27),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(27),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(27));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(30),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(30),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(30));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(31),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(31),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(31));
\GRLFPC2_0_COMB_DBGDATA_4_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(2),
dataa => N_404,
datab => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(2),
datac => \GRLFPC2_0.R.FSR.CEXC\(2));
\GRLFPC2_0_COMB_DBGDATA_4_X_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(7),
dataa => N_404,
datab => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(7),
datac => \GRLFPC2_0.R.FSR.AEXC\(2));
\GRLFPC2_0_COMB_DBGDATA_4_X_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(9),
dataa => N_404,
datab => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(9),
datac => \GRLFPC2_0.R.FSR.AEXC\(4));
\GRLFPC2_0_COMB_DBGDATA_4_X_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(3),
dataa => N_404,
datab => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(3),
datac => \GRLFPC2_0.R.FSR.CEXC\(3));
\GRLFPC2_0_COMB_DBGDATA_4_X_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(22),
dataa => N_404,
datab => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(22),
datac => \GRLFPC2_0.R.FSR.NONSTD\);
\GRLFPC2_0_WRDATA_0_X_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(54),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_392,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(54));
\GRLFPC2_0_WRDATA_0_X_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(4),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_374,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(4));
\GRLFPC2_0_WRDATA_0_X_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(29),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_399,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(29));
\GRLFPC2_0_WRDATA_0_X_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(36),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_374,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(36));
\GRLFPC2_0_WRDATA_0_X_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(61),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_399,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(61));
\GRLFPC2_0_WRDATA_0_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(1),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_371,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(1));
\GRLFPC2_0_WRDATA_0_X_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(22),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_392,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(22));
\GRLFPC2_0_WRDATA_0_X_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(33),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_371,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(33));
\GRLFPC2_0_WRDATA_0_X_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(15),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_385,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(15));
\GRLFPC2_0_WRDATA_0_X_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(18),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_388,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(18));
\GRLFPC2_0_WRDATA_0_X_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(21),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_391,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(21));
\GRLFPC2_0_WRDATA_0_X_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(47),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_385,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(47));
\GRLFPC2_0_WRDATA_0_X_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(50),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_388,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(50));
\GRLFPC2_0_WRDATA_0_X_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(53),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_391,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(53));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(29),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(29),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(29));
\GRLFPC2_0_WRDATA_0_X_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(12),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_382,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(12));
\GRLFPC2_0_WRDATA_0_X_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(24),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_394,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(24));
\GRLFPC2_0_WRDATA_0_X_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(32),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_370,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(32));
\GRLFPC2_0_WRDATA_0_X_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(44),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_382,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(44));
\GRLFPC2_0_WRDATA_0_X_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(56),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_394,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(56));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(20),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(20),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(20));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(21),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(21),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(21));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(13),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(13),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(13));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(14),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(14),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(14));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(15),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(15),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(15));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(16),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(16),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(16));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(9),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(9),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(9));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(10),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(10),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(10));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(11),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(11),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(11));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(12),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(12),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(12));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(7),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(7),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(7));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(8),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(8),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(8));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(22),
dataa => \GRLFPC2_0.COMB.V.E.STDATA2_X\,
datab => \GRLFPC2_0.R.I.INST\(22),
datac => \GRLFPC2_0.COMB.V.I.PC_1\(22));
\GRLFPC2_0_COMB_DBGDATA_4_X_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(5),
dataa => N_404,
datab => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(5),
datac => \GRLFPC2_0.R.FSR.AEXC\(0));
\GRLFPC2_0_COMB_DBGDATA_4_X_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(6),
dataa => N_404,
datab => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(6),
datac => \GRLFPC2_0.R.FSR.AEXC\(1));
\GRLFPC2_0_COMB_DBGDATA_4_X_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(8),
dataa => N_404,
datab => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(8),
datac => \GRLFPC2_0.R.FSR.AEXC\(3));
\GRLFPC2_0_WRDATA_0_X_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(5),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_375,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(5));
\GRLFPC2_0_WRDATA_0_X_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(6),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_376,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(6));
\GRLFPC2_0_WRDATA_0_X_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(37),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_375,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(37));
\GRLFPC2_0_WRDATA_0_X_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(38),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_376,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(38));
\GRLFPC2_0_COMB_DBGDATA_4_X_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(0),
dataa => N_404,
datab => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(0),
datac => \GRLFPC2_0.R.FSR.CEXC\(0));
\GRLFPC2_0_COMB_DBGDATA_4_X_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(4),
dataa => N_404,
datab => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(4),
datac => \GRLFPC2_0.R.FSR.CEXC\(4));
\GRLFPC2_0_COMB_DBGDATA_4_X_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(10),
dataa => N_404,
datab => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(10),
datac => CPO_CCZ(0));
\GRLFPC2_0_COMB_DBGDATA_4_X_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(25),
dataa => N_404,
datab => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(25),
datac => \GRLFPC2_0.R.FSR.TEM\(2));
\GRLFPC2_0_COMB_DBGDATA_4_X_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(26),
dataa => N_404,
datab => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(26),
datac => \GRLFPC2_0.R.FSR.TEM\(3));
\GRLFPC2_0_COMB_DBGDATA_4_X_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(30),
dataa => N_404,
datab => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(30),
datac => \GRLFPC2_0.R.FSR.RD\(0));
\GRLFPC2_0_COMB_DBGDATA_4_X_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(31),
dataa => N_404,
datab => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(31),
datac => \GRLFPC2_0.R.FSR.RD\(1));
\GRLFPC2_0_WRDATA_0_X_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(25),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_395,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(25));
\GRLFPC2_0_WRDATA_0_X_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(27),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_397,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(27));
\GRLFPC2_0_WRDATA_0_X_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(30),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_400,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(30));
\GRLFPC2_0_WRDATA_0_X_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(57),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_395,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(57));
\GRLFPC2_0_WRDATA_0_X_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(59),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_397,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(59));
\GRLFPC2_0_WRDATA_0_X_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(62),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_400,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(62));
\GRLFPC2_0_COMB_DBGDATA_4_X_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(23),
dataa => N_404,
datab => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(23),
datac => \GRLFPC2_0.R.FSR.TEM\(0));
\GRLFPC2_0_WRDATA_0_X_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(8),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_378,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(8));
\GRLFPC2_0_WRDATA_0_X_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(11),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_381,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(11));
\GRLFPC2_0_WRDATA_0_X_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(14),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_384,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(14));
\GRLFPC2_0_WRDATA_0_X_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(17),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_387,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(17));
\GRLFPC2_0_WRDATA_0_X_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(20),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_390,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(20));
\GRLFPC2_0_WRDATA_0_X_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(23),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_393,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(23));
\GRLFPC2_0_WRDATA_0_X_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(31),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_401,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(31));
\GRLFPC2_0_WRDATA_0_X_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(40),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_378,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(40));
\GRLFPC2_0_WRDATA_0_X_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(43),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_381,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(43));
\GRLFPC2_0_WRDATA_0_X_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(46),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_384,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(46));
\GRLFPC2_0_WRDATA_0_X_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(49),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_387,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(49));
\GRLFPC2_0_WRDATA_0_X_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(52),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_390,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(52));
\GRLFPC2_0_WRDATA_0_X_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(55),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_393,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(55));
\GRLFPC2_0_WRDATA_0_X_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(13),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_383,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(13));
\GRLFPC2_0_WRDATA_0_X_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(16),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_386,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(16));
\GRLFPC2_0_WRDATA_0_X_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(19),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_389,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(19));
\GRLFPC2_0_WRDATA_0_X_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(28),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_398,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(28));
\GRLFPC2_0_WRDATA_0_X_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(45),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_383,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(45));
\GRLFPC2_0_WRDATA_0_X_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(48),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_386,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(48));
\GRLFPC2_0_WRDATA_0_X_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(51),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_389,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(51));
\GRLFPC2_0_WRDATA_0_X_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(7),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_377,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(7));
\GRLFPC2_0_WRDATA_0_X_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(9),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_379,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(9));
\GRLFPC2_0_WRDATA_0_X_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(39),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_377,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(39));
\GRLFPC2_0_WRDATA_0_X_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(60),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_398,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(60));
\GRLFPC2_0_WRDATA_0_X_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(0),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_370,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(0));
\GRLFPC2_0_WRDATA_0_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(2),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_372,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(2));
\GRLFPC2_0_WRDATA_0_X_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(3),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_373,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(3));
\GRLFPC2_0_WRDATA_0_X_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(10),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_380,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(10));
\GRLFPC2_0_WRDATA_0_X_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(34),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_372,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(34));
\GRLFPC2_0_WRDATA_0_X_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(35),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_373,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(35));
\GRLFPC2_0_WRDATA_0_X_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.WRDATA_0_X\(42),
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => N_380,
datac => \GRLFPC2_0.COMB.WRDATA_4_X\(42));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101000011010000")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(1),
dataa => N_158,
datab => N_159,
datac => \GRLFPC2_0.R.I.INST\(1));
\GRLFPC2_0_COMB_V_E_STDATA_1_0_X_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101000011010000")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(0),
dataa => N_158,
datab => N_159,
datac => \GRLFPC2_0.R.I.INST\(0));
GRLFPC2_0_N_939_I_I_2_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC2_0.N_939_I_I_2_X\,
dataa => N_91,
datab => N_18,
datac => N_92);
GRLFPC2_0_COMB_UN1_FPCI_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC2_0.COMB.UN1_FPCI_X\,
dataa => N_368,
datab => N_367,
datac => N_18);
GRLFPC2_0_V_STATE_0_SQMUXA_1_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC2_0.V.STATE_0_SQMUXA_1_X\,
dataa => N_404,
datab => N_403,
datac => N_402);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MAPMULXFF_UN4_UNIMPMAP_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111110111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MAPMULXFF.UN4_UNIMPMAP_X\,
dataa => N_69,
datab => N_66,
datac => N_68);
GRLFPC2_0_RS1D_CNST_0_A3_0_A2_1_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC2_0.RS1D_CNST_0_A3_0_A2_1_X\,
dataa => N_68,
datab => N_67,
datac => N_66);
GRLFPC2_0_COMB_RDD_1_M14_0_A2_1_0_0_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC2_0.COMB.RDD_1.M14_0_A2_1_0_0_X\,
dataa => N_81,
datab => N_79,
datac => N_76);
GRLFPC2_0_COMB_UN1_FPCI_3_1_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC2_0.COMB.UN1_FPCI_3_1_X\,
dataa => N_159,
datab => \GRLFPC2_0.R.A.ST_RET\,
datac => \GRLFPC2_0.R.A.RS1D\);
GRLFPC2_0_COMB_UN2_HOLDN_0_A2_0_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001000")
port map (
combout => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_0_X\,
dataa => N_17,
datab => \GRLFPC2_0.R.A.MOV_RET\(15),
datac => \GRLFPC2_0.R.A.MOV_RET\(12));
\GRLFPC2_0_R_A_RF2REN_RNO_1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC2_0.COMB.V.A.RF2REN_1_0_8287_I_A4_0_0_X\,
dataa => N_89,
datab => N_90,
datac => N_79);
GRLFPC2_0_N_939_I_I_A2_0_1_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC2_0.N_939_I_I_A2_0_1_X\,
dataa => N_81,
datab => N_79,
datac => N_88);
GRLFPC2_0_R_A_LD_RNO_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC2_0.R.A.LD_0_0_G1_2_X\,
dataa => N_87,
datab => N_80,
datac => N_78);
GRLFPC2_0_COMB_ISFPOP2_1_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.ISFPOP2_1_X\,
dataa => N_352,
datab => \GRLFPC2_0.R.I.INST\(19),
datac => \GRLFPC2_0.COMB.UN1_R.I.V_0\);
GRLFPC2_0_COMB_RDD_1_M14_0_O2_0_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011100000111000")
port map (
combout => \GRLFPC2_0.COMB.RDD_1.M14_0_O2_0_X\,
dataa => N_62,
datab => N_67,
datac => N_69);
\GRLFPC2_0_COMB_V_FSR_FCC_1_0_X_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.FCC_1_0_X\(0),
dataa => N_420,
datab => \GRLFPC2_0.V.STATE_0_SQMUXA_1_X\,
datac => \GRLFPC2_0.R.I.CC\(0));
\GRLFPC2_0_COMB_V_FSR_FCC_1_0_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.FCC_1_0_X\(1),
dataa => N_421,
datab => \GRLFPC2_0.V.STATE_0_SQMUXA_1_X\,
datac => \GRLFPC2_0.R.I.CC\(1));
\GRLFPC2_0_RS1_1_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => RFI2_RD1ADDRZ(0),
dataa => N_402,
datab => N_406,
datac => \GRLFPC2_0.COMB.RS1_1\(1));
\GRLFPC2_0_RS1_1_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => RFI2_RD1ADDRZ(1),
dataa => N_402,
datab => N_407,
datac => \GRLFPC2_0.COMB.RS1_1\(2));
\GRLFPC2_0_RS1_1_X_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => RFI2_RD1ADDRZ(2),
dataa => N_402,
datab => N_408,
datac => \GRLFPC2_0.COMB.RS1_1\(3));
\GRLFPC2_0_RS1_1_X_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => RFI2_RD1ADDRZ(3),
dataa => N_402,
datab => N_409,
datac => \GRLFPC2_0.COMB.RS1_1\(4));
\GRLFPC2_0_RS2_1_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => RFI2_RD2ADDRZ(0),
dataa => N_402,
datab => N_406,
datac => \GRLFPC2_0.COMB.RS2_1\(1));
\GRLFPC2_0_RS2_1_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => RFI2_RD2ADDRZ(1),
dataa => N_402,
datab => N_407,
datac => \GRLFPC2_0.COMB.RS2_1\(2));
\GRLFPC2_0_RS2_1_X_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => RFI2_RD2ADDRZ(2),
dataa => N_402,
datab => N_408,
datac => \GRLFPC2_0.COMB.RS2_1\(3));
\GRLFPC2_0_RS2_1_X_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => RFI2_RD2ADDRZ(3),
dataa => N_402,
datab => N_409,
datac => \GRLFPC2_0.COMB.RS2_1\(4));
GRLFPC2_0_WRADDR_0_SQMUXA_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
dataa => \GRLFPC2_0.COMB.UN1_FPCI_X\,
datab => \GRLFPC2_0.R.X.AFSR\,
datac => \GRLFPC2_0.R.X.LD\);
GRLFPC2_0_R_X_AFSR_RNIOEMG: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC2_0.V.FSR.NONSTD_0_SQMUXA_6_X\,
dataa => \GRLFPC2_0.COMB.UN1_FPCI_X\,
datab => \GRLFPC2_0.R.X.AFSR\,
datac => \GRLFPC2_0.R.X.LD\);
\GRLFPC2_0_COMB_V_I_RES_6_X_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001000010010")
port map (
combout => \GRLFPC2_0.COMB.V.I.RES_6_X\(63),
dataa => N_133,
datab => N_134,
datac => \GRLFPC2_0.FPI.OP2_X\(63));
GRLFPC2_0_COMB_V_I_EXEC_4_IV_0_A2_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000010110000")
port map (
combout => \GRLFPC2_0.COMB.V.I.EXEC_4_IV_0_A2_X\,
dataa => \GRLFPC2_0.COMB.UN1_FPCI_X\,
datab => \GRLFPC2_0.R.X.SEQERR\,
datac => \GRLFPC2_0.R.I.EXEC\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MAPMULXFF_UNIMPMAP_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001000010010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MAPMULXFF.UNIMPMAP_X\,
dataa => N_76,
datab => N_70,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MAPMULXFF.UN4_UNIMPMAP_X\);
GRLFPC2_0_RS1V_0_SQMUXA_0_A2_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001000010010000")
port map (
combout => \GRLFPC2_0.RS1V_0_SQMUXA_0_A2_X\,
dataa => N_76,
datab => N_77,
datac => \GRLFPC2_0.R.A.ST_RET_0_0_G1\);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_2_A_X_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011101000111")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_2_A_X\(0),
dataa => N_410,
datab => \GRLFPC2_0.V.STATE_0_SQMUXA_1_X\,
datac => \GRLFPC2_0.R.I.EXC\(0));
\GRLFPC2_0_COMB_V_FSR_CEXC_1_2_A_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011101000111")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_2_A_X\(2),
dataa => N_412,
datab => \GRLFPC2_0.V.STATE_0_SQMUXA_1_X\,
datac => \GRLFPC2_0.R.I.EXC\(2));
\GRLFPC2_0_COMB_V_FSR_CEXC_1_2_A_X_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011101000111")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_2_A_X\(4),
dataa => N_414,
datab => \GRLFPC2_0.V.STATE_0_SQMUXA_1_X\,
datac => \GRLFPC2_0.R.I.EXC\(4));
\GRLFPC2_0_COMB_V_FSR_CEXC_1_2_A_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011101000111")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_2_A_X\(1),
dataa => N_411,
datab => \GRLFPC2_0.V.STATE_0_SQMUXA_1_X\,
datac => \GRLFPC2_0.R.I.EXC\(1));
\GRLFPC2_0_COMB_V_FSR_CEXC_1_2_A_X_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011101000111")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_2_A_X\(3),
dataa => N_413,
datab => \GRLFPC2_0.V.STATE_0_SQMUXA_1_X\,
datac => \GRLFPC2_0.R.I.EXC\(3));
GRLFPC2_0_V_STATE_1_SQMUXA_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100110001001100")
port map (
combout => \GRLFPC2_0.V.STATE_1_SQMUXA_X\,
dataa => N_438,
datab => N_8,
datac => \GRLFPC2_0.V.STATE_0_SQMUXA_1_X\);
GRLFPC2_0_COMB_RDD_1_M14_0_A2_1_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC2_0.COMB.RDD_1.M14_0_A2_1_X\,
dataa => N_77,
datab => \GRLFPC2_0.COMB.RDD_1.M14_0_A2_1_0_0_X\,
datac => \GRLFPC2_0.COMB.RDD_1.M14_0_A2_1_1\);
GRLFPC2_0_R_X_SEQERR_RNI85A8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000101010001010")
port map (
combout => \GRLFPC2_0.R.I.V_1_0_G2_0_0_X\,
dataa => N_8,
datab => \GRLFPC2_0.COMB.UN1_FPCI_X\,
datac => \GRLFPC2_0.R.X.SEQERR\);
GRLFPC2_0_FPI_LDOP_0_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110111111101")
port map (
combout => \GRLFPC2_0.FPI.LDOP_0_X\,
dataa => N_8,
datab => \GRLFPC2_0.R.MK.RST2\,
datac => \GRLFPC2_0.COMB.V.MK.RST_1_0_A2\);
GRLFPC2_0_R_MK_BUSY2_RET_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.R.MK.BUSY2_RET_0_0_A2_0_G0_X\,
dataa => N_8,
datab => \GRLFPC2_0.COMB.ANNULFPU_1_U_0_O2\);
\GRLFPC2_0_R_A_RF2REN_RNO_0_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC2_0.COMB.V.A.RF2REN_1_0_8287_I_A4_0_X\,
dataa => N_81,
datab => \GRLFPC2_0.COMB.V.A.RF2REN_1_0_8287_I_A4_0_0_X\,
datac => \GRLFPC2_0.N_939_I_I_O2\);
\GRLFPC2_0_R_FSR_FTT_RNO_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC2_0.R.FSR.FTT_0_0_2__G1_X\,
dataa => N_8,
datab => \GRLFPC2_0.R.FSR.FTT_0_0_2__G1_A\,
datac => \GRLFPC2_0.N_1570_I_I_A2\);
GRLFPC2_0_COMB_RS2D_1_IV_0_O2_RNIKKJ6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.R.A.RS2D_0_0_G1_0_X\,
dataa => N_70,
datab => \GRLFPC2_0.COMB.RS2D_1_IV_0_O2\);
GRLFPC2_0_V_FSR_AEXC_1_SQMUXA_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000100")
port map (
combout => \GRLFPC2_0.V.FSR.AEXC_1_SQMUXA_X\,
dataa => \GRLFPC2_0.V.STATE_0_SQMUXA_1_X\,
datab => \GRLFPC2_0.V.FSR.NONSTD_0_SQMUXA_6_X\,
datac => \GRLFPC2_0.COMB.V.FSR.FCC8\);
GRLFPC2_0_COMB_UN7_RS2V_0_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC2_0.COMB.UN7_RS2V_0_X\,
dataa => \GRLFPC2_0.R.A.RS2D_0_0_G1\,
datab => \GRLFPC2_0.COMB.RS2_1\(0));
GRLFPC2_0_V_FSR_AEXC_2_SQMUXA_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA_X\,
dataa => \GRLFPC2_0.V.STATE_0_SQMUXA_1_X\,
datab => \GRLFPC2_0.V.FSR.NONSTD_0_SQMUXA_6_X\,
datac => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA_1\);
\GRLFPC2_0_COMB_RF1REN_1_0_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.RF1REN_1_0_X\(1),
dataa => N_17,
datab => \GRLFPC2_0.R.A.RF1REN\(1),
datac => \GRLFPC2_0.COMB.V.A.RF1REN_1\(1));
\GRLFPC2_0_COMB_RF2REN_1_0_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.COMB.RF2REN_1_0_X\(1),
dataa => N_17,
datab => \GRLFPC2_0.R.A.RF2REN\(1),
datac => \GRLFPC2_0.COMB.V.A.RF2REN_1\(1));
GRLFPC2_0_COMB_WREN1_10_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010100010101000")
port map (
combout => \GRLFPC2_0.COMB.WREN1_10_X\,
dataa => N_17,
datab => \GRLFPC2_0.COMB.WREN1_9_IV_0\,
datac => \GRLFPC2_0.COMB.WREN1_9_IV_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000010000001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW_0_0_7__G0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_IV\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW_0_0_7__G1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_IV\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110111111101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CONDMUXMULXFF.UN4_NOTSQRTLFTCC\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA_RNIF9664: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_58__G0\,
dataa => \GRLFPC2_0.FPI.LDOP_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_317__G1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_58__G2_M9_I_M4\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_RNIRFK3_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000001010000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_0_0_3__G0_I\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_IV\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_27: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111011110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN7_FEEDBACK_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_24\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27_D_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_0_0_13__G0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12),
datab => NN_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_I_M_3950\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_0_0_13__G0_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_2_IV_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_IV\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_AREGSIGN_SEL_INV\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_IV_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_I_M\(13));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD55_RNIQGGR1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000110011111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_58__G2_M9_I_M4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD55\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_58__G2_M9_I_M4_A\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD57_RNIRC6F1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_58__G2_M9_I_M4_A\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD57\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_58__G2TT_M2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_27_D_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111011110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27_D_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(49),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_21\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27_D\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_0_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000101011001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_0_0_13__G0_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(13),
datab => \GRLFPC2_0.FPI.OP1_X\(63),
datac => \GRLFPC2_0.FPI.LDOP_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_AREGSIGN_SEL_INV_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_1_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_59__G0_XX\,
dataa => \GRLFPC2_0.FPI.LDOP_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_318__G1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(59));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_27_D: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_27_D\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(49),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_15\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_18\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4_A\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_A_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4_A\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_2_IV_RNO_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_I_M\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(22),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SFTLFT.UN4_TEMP\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_I_M_3950\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN28_STKOUT_RNIGO5K6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN22_NOTPROP_0_S\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1_5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN28_STKOUT\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_UN4_XZBREGLOADEN_RNIN2P11: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111101110111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_58__G2TT_M2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLBREGXZ.UN4_XZBREGLOADEN\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.WQSCTRL_0\(67),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SS0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111000010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLBREGXZ.UN4_XZBREGLOADEN\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.WQSCTRL_0\(67),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_24: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110011011100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_24\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN30_CONDITIONAL_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_18: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110100100001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_18\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_17\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_2_IV_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110000001101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_IV_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(0),
datab => \GRLFPC2_0.FPI.OP2_X\(63),
datac => \GRLFPC2_0.FPI.LDOP_REP5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_IV_0_A\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_2_IV_0_A_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_IV_0_A\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(22),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.SIGNRESULT\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.WQSCTRL_0_3947\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_316_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_316__G1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_114_C0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_0\(56));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_1_RNIVD872: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_317__G1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_114_C0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_0\(56));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_1_RNIMN8B2_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_318__G1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_114_SUM0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_116_C0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_3_RNI3VCR2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_319__G1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_60_C1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_116_SUM0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2S2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.WQSCTRL_0_3947\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_50_1.SUM_0\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_1.SUM_0\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_AREGSIGN_SEL_INV_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001111111111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_AREGSIGN_SEL_INV_1\,
dataa => NN_2,
datab => \GRLFPC2_0.FPI.LDOP_REP5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.WQSCTRL_0_3947\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_AREGSIGN_SEL_INV: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000111111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_AREGSIGN_SEL_INV\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(22),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SFTLFT.UN4_TEMP\,
datac => \GRLFPC2_0.FPI.LDOP_REP5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.WQSCTRL_0\(67));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_REP4_RNIOF0I: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_I_M_3950\,
dataa => \GRLFPC2_0.FPI.LDOP_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.WQSCTRL_0_3947\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLAREGXZ.UN5_XZAREGLOADEN_0\,
datac => \GRLFPC2_0.FPI.LDOP_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.WQSCTRL_0\(67));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN2_MIXOIN_3_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100110011101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_3\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN22_NOTPROP_0_S\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.GEN_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_SUM4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_2\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN28_STKOUT: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101101011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN28_STKOUT\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN22_NOTPROP_0_S\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN36_STKGEN_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_SUM4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_2\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_12_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G_32\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN20_STKOUT_RNIUQTT3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1_5\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN16_NOTPROP_0_S\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_1\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN20_STKOUT\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_51\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_50\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_53\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_55\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN30_CONDITIONAL_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN30_CONDITIONAL_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN30_CONDITIONAL_0_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN30_CONDITIONAL_M5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_1_SQMUXA_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLBREGXZ.UN4_XZBREGLOADEN\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLBREGXZ.XZBREGLC_2\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.WQSCTRL_0_3947\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23_1_SUM_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011101111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_1.SUM_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_114_C0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_0\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_50_1_SUM_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011101111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_50_1.SUM_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_114_C0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_0\(56));
GRLFPC2_0_COMB_WREN1_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111100100000")
port map (
combout => RFI1_WRENZ,
dataa => N_402,
datab => N_405,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.COMB.WREN1_10_X\);
GRLFPC2_0_COMB_WREN2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRENZ,
dataa => N_402,
datab => N_405,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.COMB.WREN2_10\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_261__G0_I_X4_0_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_262__G0_I_X4_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_258_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011101111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_258__G0_I_X4_0_0_0_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_114_C0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_0\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_RNI8CAG_68_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111000000110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.WQSCTRL_0\(67),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.WQSCTRL\(68),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD57\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_GEN_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000111100001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.GEN_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.GEN_3_A\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_ADD2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_GEN_3_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100110011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.GEN_3_A\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_C1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_ADD1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_55: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_55\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_35\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_36\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_45\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_46\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001100")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV\(4),
dataa => \GRLFPC2_0.R.FSR.AEXC\(4),
datab => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV_0\(4),
datac => \GRLFPC2_0.COMB.V.FSR.AEXC_6_I_M\(4),
datad => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA_X\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001100")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV\(0),
dataa => \GRLFPC2_0.R.FSR.AEXC\(0),
datab => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV_0\(0),
datac => \GRLFPC2_0.COMB.V.FSR.AEXC_6_I_M\(0),
datad => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA_X\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001100")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV\(1),
dataa => \GRLFPC2_0.R.FSR.AEXC\(1),
datab => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV_0\(1),
datac => \GRLFPC2_0.COMB.V.FSR.AEXC_6_I_M\(1),
datad => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA_X\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001100")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV\(2),
dataa => \GRLFPC2_0.R.FSR.AEXC\(2),
datab => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV_0\(2),
datac => \GRLFPC2_0.COMB.V.FSR.AEXC_6_I_M\(2),
datad => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA_X\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001100")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV\(3),
dataa => \GRLFPC2_0.R.FSR.AEXC\(3),
datab => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV_0\(3),
datac => \GRLFPC2_0.COMB.V.FSR.AEXC_6_I_M\(3),
datad => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA_X\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_3_RNI3VCR2_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011101111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_262__G0_I_X4_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_60_C1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_116_SUM0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_1_RNIMN8B2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011101111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_261__G0_I_X4_0_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_114_SUM0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_116_C0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN36_STKGEN_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111010000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN36_STKGEN_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_C1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_ADD1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_ADD2\);
GRLFPC2_0_COMB_WREN2_10: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101000")
port map (
combout => \GRLFPC2_0.COMB.WREN2_10\,
dataa => N_17,
datab => \GRLFPC2_0.COMB.WREN2_9_IV_0\,
datac => \GRLFPC2_0.WREN1_0_SQMUXA_1\,
datad => \GRLFPC2_0.COMB.WRADDR_5_M\(0));
\GRLFPC2_0_COMB_RF1REN_1_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111110110000")
port map (
combout => RFI1_REN1Z,
dataa => N_404,
datab => N_403,
datac => N_402,
datad => \GRLFPC2_0.COMB.RF1REN_1_0_X\(1));
\GRLFPC2_0_COMB_RF1REN_1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111110110000")
port map (
combout => RFI1_REN2Z,
dataa => N_404,
datab => N_403,
datac => N_402,
datad => \GRLFPC2_0.COMB.RF1REN_1_0_0\(2));
\GRLFPC2_0_COMB_RF2REN_1_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111110110000")
port map (
combout => RFI2_REN1Z,
dataa => N_404,
datab => N_403,
datac => N_402,
datad => \GRLFPC2_0.COMB.RF2REN_1_0_X\(1));
\GRLFPC2_0_COMB_RF2REN_1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111110110000")
port map (
combout => RFI2_REN2Z,
dataa => N_404,
datab => N_403,
datac => N_402,
datad => \GRLFPC2_0.COMB.RF2REN_1_0\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_RNIJ1P9_68_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111001101110011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.WQSCTRL_0_3947\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.WQSCTRL\(68),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD57\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_RNIIVV94: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001011111101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_SUM4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_C1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_ADD1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_ADD2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN20_STKOUT: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101101011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN20_STKOUT\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN16_NOTPROP_0_S\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN27_STKGEN_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_SUM3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_RESULT_U_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100111011000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_U\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(49),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G_31_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_0\(1));
\GRLFPC2_0_R_A_RF1REN_RNO_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001001100")
port map (
combout => \GRLFPC2_0.COMB.V.A.RF1REN_1_8259_I\,
dataa => \GRLFPC2_0.COMB.V.A.RF1REN_1_8259_I_A5_0\,
datab => \GRLFPC2_0.COMB.V.A.RF1REN_1_8259_I_0\,
datac => \GRLFPC2_0.COMB.RS1_1_0_X\(0),
datad => \GRLFPC2_0.N_939_I_I_A2\);
\GRLFPC2_0_R_A_RF2REN_RNO_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011000100")
port map (
combout => \GRLFPC2_0.COMB.V.A.RF2REN_1_8311_I\,
dataa => \GRLFPC2_0.COMB.V.A.RF1REN_1_8259_I_A5_0\,
datab => \GRLFPC2_0.COMB.V.A.RF2REN_1_8311_I_0\,
datac => \GRLFPC2_0.COMB.RS1_1_0_X\(0),
datad => \GRLFPC2_0.N_939_I_I_A2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_3_RNI6HOV: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_114_C0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_58_C0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58_0\(56));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_3_RNICO8J1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_60_C1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_58_SUM0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_60_C0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_3_RNIBHC41_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_116_C0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_58_C0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58_0\(56));
\GRLFPC2_0_COMB_RF1REN_1_0_0_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111010001000100")
port map (
combout => \GRLFPC2_0.COMB.RF1REN_1_0_0\(2),
dataa => N_17,
datab => \GRLFPC2_0.R.A.RF1REN\(2),
datac => \GRLFPC2_0.COMB.RF1REN_1_0_0_A2_1\(2),
datad => \GRLFPC2_0.COMB.FPOP_0_0_O2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(173),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datac => \GRLFPC2_0.FPI.LDOP_REP5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN2_MIXOIN_2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000011110111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_2\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN16_NOTPROP_0_S\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_SUM3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.GEN_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_RESULT_0_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111011110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_0\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN7_FEEDBACK_0_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN7_FEEDBACK_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SFTLFT.AREGXORBREG_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.REEXCOVUV.UN3_LOCUV\);
\GRLFPC2_0_COMB_RF2REN_1_0_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010011100100")
port map (
combout => \GRLFPC2_0.COMB.RF2REN_1_0\(2),
dataa => N_17,
datab => \GRLFPC2_0.R.A.RF2REN\(2),
datac => \GRLFPC2_0.COMB.UN7_RS2V_0_X\,
datad => \GRLFPC2_0.N_939_I_I_A2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_21: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001001110011100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_21\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN30_CONDITIONAL_0_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN30_CONDITIONAL_0_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD11\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD12\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN12_STKOUT_RNID9352: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN10_NOTPROP_0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN12_STKOUT\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_46: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_46\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(30),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_8\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_13\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_45: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_45\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_5\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_6\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN18_XZXBUS_18_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_33\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_0_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110010101111")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV_0\(3),
dataa => N_418,
datab => N_378,
datac => \GRLFPC2_0.V.STATE_0_SQMUXA_1_X\,
datad => \GRLFPC2_0.V.FSR.AEXC_1_SQMUXA_X\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110010101111")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV_0\(0),
dataa => N_415,
datab => N_375,
datac => \GRLFPC2_0.V.STATE_0_SQMUXA_1_X\,
datad => \GRLFPC2_0.V.FSR.AEXC_1_SQMUXA_X\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_0_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110010101111")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV_0\(4),
dataa => N_419,
datab => N_379,
datac => \GRLFPC2_0.V.STATE_0_SQMUXA_1_X\,
datad => \GRLFPC2_0.V.FSR.AEXC_1_SQMUXA_X\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_0_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110010101111")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV_0\(1),
dataa => N_416,
datab => N_376,
datac => \GRLFPC2_0.V.STATE_0_SQMUXA_1_X\,
datad => \GRLFPC2_0.V.FSR.AEXC_1_SQMUXA_X\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_0_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110010101111")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV_0\(2),
dataa => N_417,
datab => N_377,
datac => \GRLFPC2_0.V.STATE_0_SQMUXA_1_X\,
datad => \GRLFPC2_0.V.FSR.AEXC_1_SQMUXA_X\);
GRLFPC2_0_COMB_WREN1_9_IV_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111010011110100")
port map (
combout => \GRLFPC2_0.COMB.WREN1_9_IV_1\,
dataa => \GRLFPC2_0.COMB.WRADDR_5_X\(0),
datab => \GRLFPC2_0.WREN1_1_SQMUXA_2\,
datac => \GRLFPC2_0.WREN1_0_SQMUXA_1\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_RNO_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_6_I_M\(4),
dataa => \GRLFPC2_0.V.STATE_0_SQMUXA_1_X\,
datab => \GRLFPC2_0.R.FSR.AEXC\(4),
datac => \GRLFPC2_0.R.I.EXC\(4),
datad => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA_1\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_RNO_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_6_I_M\(2),
dataa => \GRLFPC2_0.V.STATE_0_SQMUXA_1_X\,
datab => \GRLFPC2_0.R.FSR.AEXC\(2),
datac => \GRLFPC2_0.R.I.EXC\(2),
datad => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA_1\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_RNO_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_6_I_M\(1),
dataa => \GRLFPC2_0.V.STATE_0_SQMUXA_1_X\,
datab => \GRLFPC2_0.R.FSR.AEXC\(1),
datac => \GRLFPC2_0.R.I.EXC\(1),
datad => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA_1\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_RNO_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_6_I_M\(0),
dataa => \GRLFPC2_0.V.STATE_0_SQMUXA_1_X\,
datab => \GRLFPC2_0.R.FSR.AEXC\(0),
datac => \GRLFPC2_0.R.I.EXC\(0),
datad => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA_1\);
\GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_RNO_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.AEXC_6_I_M\(3),
dataa => \GRLFPC2_0.V.STATE_0_SQMUXA_1_X\,
datab => \GRLFPC2_0.R.FSR.AEXC\(3),
datac => \GRLFPC2_0.R.I.EXC\(3),
datad => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA_1\);
\GRLFPC2_0_R_A_RF2REN_RNO_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010001100")
port map (
combout => \GRLFPC2_0.COMB.V.A.RF2REN_1_0_8287_I\,
dataa => N_57,
datab => \GRLFPC2_0.COMB.RS1_1_SN_M2_I_A2\,
datac => \GRLFPC2_0.COMB.V.A.RF2REN_1_0_8287_I_O4_0\,
datad => \GRLFPC2_0.COMB.V.A.RF2REN_1_0_8287_I_A4_0_X\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_3_RNI6HOV_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011101111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_114_SUM0_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_58_C0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58_0\(56));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2_2_RNIP70T: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011101111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_0\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_58_C0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58_0\(56));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_3_RNIBHC41: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011101111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_116_SUM0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_58_C0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58_0\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(115),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(57));
\GRLFPC2_0_COMB_V_A_RF1REN_1_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010001100")
port map (
combout => \GRLFPC2_0.COMB.V.A.RF1REN_1\(1),
dataa => \GRLFPC2_0.COMB.RS1D_1_U\,
datab => \GRLFPC2_0.COMB.RS1V_1_IV\,
datac => \GRLFPC2_0.COMB.RS1_1\(0),
datad => \GRLFPC2_0.N_939_I_I_A2\);
\GRLFPC2_0_COMB_V_A_RF2REN_1_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011001000")
port map (
combout => \GRLFPC2_0.COMB.V.A.RF2REN_1\(1),
dataa => \GRLFPC2_0.COMB.RS1D_1_U\,
datab => \GRLFPC2_0.COMB.RS1V_1_IV\,
datac => \GRLFPC2_0.COMB.RS1_1\(0),
datad => \GRLFPC2_0.N_939_I_I_A2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_RNI3IOA2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110100110010110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN22_NOTPROP_0_S\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_C1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_ADD1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_GEN_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100011111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.GEN_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_SUM1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_C1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN19_GEN\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN3_LOCUV: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110111011101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.REEXCOVUV.UN3_LOCUV\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD12\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_13: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_13\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_7\);
\GRLFPC2_0_R_A_RF1REN_RNO_0_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111011100000000")
port map (
combout => \GRLFPC2_0.COMB.V.A.RF1REN_1_8259_I_0\,
dataa => N_82,
datab => \GRLFPC2_0.RS1V_0_SQMUXA_0_A2_X\,
datac => \GRLFPC2_0.RS1D_CNST_0_A2\,
datad => \GRLFPC2_0.COMB.RS1V_1_IV\);
\GRLFPC2_0_R_A_RF2REN_RNO_0_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111000000000")
port map (
combout => \GRLFPC2_0.COMB.V.A.RF2REN_1_8311_I_0\,
dataa => \GRLFPC2_0.COMB.RS1_1_SN_M2_I_A2\,
datab => \GRLFPC2_0.COMB.RS1_1_1_X\(0),
datac => \GRLFPC2_0.RS1D_CNST_0_A2\,
datad => \GRLFPC2_0.COMB.RS1V_1_IV\);
\GRLFPC2_0_COMB_RF1REN_1_0_0_A2_1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100010001000")
port map (
combout => \GRLFPC2_0.COMB.RF1REN_1_0_0_A2_1\(2),
dataa => \GRLFPC2_0.COMB.RS1_1_SN_M2_I_A2\,
datab => N_17,
datac => \GRLFPC2_0.COMB.V.A.RF2REN_1_0_8287_I_O4_0\,
datad => \GRLFPC2_0.COMB.RS2_1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_3_RNICO8J1_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011101111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_60_SUM1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_58_SUM0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_60_C0\);
GRLFPC2_0_V_FSR_CEXC_3_SQMUXA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC2_0.V.FSR.CEXC_3_SQMUXA\,
dataa => \GRLFPC2_0.V.STATE_0_SQMUXA_1_X\,
datab => \GRLFPC2_0.V.FSR.NONSTD_0_SQMUXA_6_X\,
datac => \GRLFPC2_0.N_1570_I_I_A2\,
datad => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_NE: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_8\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_9\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN19_GEN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN19_GEN\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_C0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_SUM1_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN20_GEN\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN27_STKGEN_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111010000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN27_STKGEN_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_SUM0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_C0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_SUM1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.STARTSHFT.UN3_NOTRESETORUNIMP\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW\(77),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.STARTSHFT.UN3_NOTRESETORUNIMP\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_BUSYMULXFF_UN2_TEMP: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111111111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.BUSYMULXFF.UN2_TEMP\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW\(77),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.BUSYMULXFF.UN2_TEMP_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28\);
GRLFPC2_0_R_I_EXEC_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.R.I.EXEC_0_0_G1\,
dataa => \GRLFPC2_0.R.I.V_1_0_G2_0\,
datab => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2\,
datac => \GRLFPC2_0.COMB.V.I.EXEC\,
datad => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA_1\);
GRLFPC2_0_R_I_V_RNO_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110111111111")
port map (
combout => \GRLFPC2_0.R.I.V_1_0_G0_I_O4\,
dataa => \GRLFPC2_0.R.I.V_1_0_G2_0\,
datab => \GRLFPC2_0.N_1570_I_I_A2\,
datac => G_8482,
datad => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA_1\);
GRLFPC2_0_V_FSR_AEXC_1_SQMUXA_0_RNIJS9I1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011111101")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_SN_M3\,
dataa => \GRLFPC2_0.V.FSR.AEXC_1_SQMUXA_0\,
datab => \GRLFPC2_0.N_1570_I_I_A2\,
datac => \GRLFPC2_0.COMB.V.FSR.FCC8\,
datad => \GRLFPC2_0.V.FSR.CEXC_3_SQMUXA\);
GRLFPC2_0_COMB_WREN2_10_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.COMB.WRADDR_5_M\(0),
dataa => \GRLFPC2_0.COMB.WRADDR_5_X\(0),
datab => \GRLFPC2_0.WREN1_1_SQMUXA_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000110100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_0\);
\GRLFPC2_0_R_FSR_FCC_RNO_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110011011000")
port map (
combout => \GRLFPC2_0.R.FSR.FCC_0_0_0__G1\,
dataa => \GRLFPC2_0.V.STATE_0_SQMUXA_1_X\,
datab => \GRLFPC2_0.COMB.V.FSR.FCC_1_0_X\(0),
datac => \GRLFPC2_0.COMB.V.FSR.FCC_1_1_X\(0),
datad => \GRLFPC2_0.COMB.V.FSR.FCC8\);
\GRLFPC2_0_R_FSR_FCC_RNO_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110011011000")
port map (
combout => \GRLFPC2_0.R.FSR.FCC_0_0_1__G1\,
dataa => \GRLFPC2_0.V.STATE_0_SQMUXA_1_X\,
datab => \GRLFPC2_0.COMB.V.FSR.FCC_1_0_X\(1),
datac => \GRLFPC2_0.COMB.V.FSR.FCC_1_1_X\(1),
datad => \GRLFPC2_0.COMB.V.FSR.FCC8\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN12_STKOUT: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111011100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN12_STKOUT\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN18_STKGEN_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN10_NOTPROP_0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.NOTPROP_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_3_RNILB2R1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001011111101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_SUM3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_SUM0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_C0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_SUM1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN2_MIXOIN_1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011101000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.GEN_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.NOTPROP_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_53: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_53\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_37\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_38\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_49\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_8\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111101101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_8\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_6\);
\GRLFPC2_0_R_I_EXC_RNO_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.R.I.EXC_2_0_2__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(38),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(40),
datad => \GRLFPC2_0.R.I.EXC_0\(0));
GRLFPC2_0_COMB_RS2D_1_IV_0_O2_RNIJTLO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.R.A.RS2D_0_0_G1\,
dataa => N_63,
datab => N_62,
datac => \GRLFPC2_0.COMB.RS1_1_SN_M2_I_A2\,
datad => \GRLFPC2_0.R.A.RS2D_0_0_G1_0_X\);
GRLFPC2_0_COMB_FPDECODE_RS1D5_0_A2_RNIJBPT: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100001001100")
port map (
combout => \GRLFPC2_0.COMB.V.A.RF1REN_1_8259_I_A5_0\,
dataa => N_76,
datab => \GRLFPC2_0.COMB.RS1_1_SN_M2_I_A2\,
datac => \GRLFPC2_0.COMB.FPDECODE.RS1D5_0_A2\,
datad => \GRLFPC2_0.RS1D_CNST_0_A2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_1_C: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_C\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.UN4_TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.TEMP_25\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.STARTSHFT.UN3_NOTRESETORUNIMP\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_PCTRL_NEW_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW\(77),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.UN3_TEMP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.STARTSHFT.UN3_NOTRESETORUNIMP\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_RNIO4M01_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_C1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_C0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_ADD0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_RNIOTCP: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_58_C0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_2_C0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_RNIFKJL: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_60_C0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_2_C0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1_0\);
GRLFPC2_0_COMB_WREN125_1_RNIB8Q81: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC2_0.WREN1_0_SQMUXA_1\,
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.COMB.V.STATE\,
datac => \GRLFPC2_0.COMB.V.STATE_7_IV_I\(0),
datad => \GRLFPC2_0.COMB.WREN125_1\);
GRLFPC2_0_WREN1_1_SQMUXA_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC2_0.WREN1_1_SQMUXA_2\,
dataa => \GRLFPC2_0.COMB.RDD_2\,
datab => \GRLFPC2_0.COMB.V.STATE\,
datac => \GRLFPC2_0.COMB.V.STATE_7_IV_I\(0),
datad => \GRLFPC2_0.COMB.WREN125_1\);
GRLFPC2_0_V_FSR_AEXC_2_SQMUXA_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011101111")
port map (
combout => \GRLFPC2_0.V.FSR.AEXC_2_SQMUXA_1\,
dataa => \GRLFPC2_0.COMB.V.STATE\,
datab => \GRLFPC2_0.COMB.V.STATE_7_IV_I\(0),
datac => \GRLFPC2_0.COMB.WREN125_1\,
datad => \GRLFPC2_0.COMB.V.FSR.FCC8\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(171),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datac => \GRLFPC2_0.FPI.LDOP_REP5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(45),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(45),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(46),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(46),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(23),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(22),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(16),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(14),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(14));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(41),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(24),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(25));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(12),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(10),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(21),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(21),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(26),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(50),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(50));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(39),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(43),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(37),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(28),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(35),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(35));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(20),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(20));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(30),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(15),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(40),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(40),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(40));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(172),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datac => \GRLFPC2_0.FPI.LDOP_REP5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(47));
GRLFPC2_0_R_E_SEQERR_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111100001000")
port map (
combout => \GRLFPC2_0.R.E.SEQERR_0_0_G1\,
dataa => \GRLFPC2_0.COMB.SEQERR.UN3_QNE_2\,
datab => \GRLFPC2_0.COMB.SEQERR.UN3_QNE_3\,
datac => \GRLFPC2_0.COMB.UN4_LOCK_0\,
datad => \GRLFPC2_0.COMB.SEQERR.SEQERR_0_A3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN20_GEN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN20_GEN\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_SUM0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_C0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_SUM1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_GEN_2_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_C1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_SUM0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_C0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_GEN_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.GEN_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP_1_SUM0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP_1_C0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_SUM0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(38));
GRLFPC2_0_COMB_RS1V_1_IV: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111100000")
port map (
combout => \GRLFPC2_0.COMB.RS1V_1_IV\,
dataa => N_89,
datab => N_90,
datac => \GRLFPC2_0.RS1V_0_SQMUXA_0_A2_X\,
datad => \GRLFPC2_0.UN1_FPOP7_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_15: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_15\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_14\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_7\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(19));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_BUSYMULXFF_UN2_TEMP_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.BUSYMULXFF.UN2_TEMP_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(68),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(70),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.UN3_TEMP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.STARTSHFT.UN2_NOTDECODEDUNIMP\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_43_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(66),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.STARTSHFT.UN3_NOTDECODEDUNIMP\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_51: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_51\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_31\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_32\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_29\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_30\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_50: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_50\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_42\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_41\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_49: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_49\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_21\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_24\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_23\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_22\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_35: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_35\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN18_XZXBUS_13_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_12\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001001001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_5\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(7));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001001001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001001001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(10),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000110000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_3_M4_I_X2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(0));
GRLFPC2_0_COMB_V_FSR_FCC8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.FCC8\,
dataa => \GRLFPC2_0.R.I.V\,
datab => \GRLFPC2_0.COMB.ISFPOP2_1_X\,
datac => \GRLFPC2_0.COMB.V.I.EXEC\,
datad => \GRLFPC2_0.COMB.UN1_V.STATE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_65_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100111111101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW_2_0_65__G0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(66),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(64),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(68),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.STARTSHFT.UN3_NOTDECODEDUNIMP\);
GRLFPC2_0_COMB_RS2D_1_IV_0_O2_RNIBTB8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110111111111")
port map (
combout => \GRLFPC2_0.COMB.V.A.RF2REN_1_0_8287_I_O4_0\,
dataa => N_63,
datab => N_62,
datac => N_70,
datad => \GRLFPC2_0.COMB.RS2D_1_IV_0_O2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_0_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_4\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_13\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_18\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_23\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_19\(47),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_21\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_18\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_20\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_1_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_8\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_9\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_14\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_19\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_20\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_22\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_21\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_23\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_16\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_20\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_17\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_22\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_17\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_18\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_19\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_A\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_A\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_8645\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_16\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_6\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_14\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_10\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_9\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_18\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_22\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_18\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_19\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_23\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_10\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_11\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_14\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_16\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_40__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_3_I_O2\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_12_0_A2\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_0\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_39__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_1\(38),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_39__G2_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_0\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2\(38));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_9\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_12\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_8\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_14\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_8\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_9\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_12\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_14\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_12\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_13\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_19\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_20\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_7\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_11\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_20_4_RNI2RVV9_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_16\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_17\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_24\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_23\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_2_RNI808A3_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_6\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_10\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_8\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_RNIBLKR_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_16__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_16__G2_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1162\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_4\(50),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2\(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_RNIOTCP_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011101111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_58_SUM0_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_2_C0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_58_0_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011101111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.SI_58_0\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_2_C0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1_0\);
\GRLFPC2_0_R_I_EXC_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000110000001110")
port map (
combout => \GRLFPC2_0.R.I.EXC_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN11_INEXACT_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN2_INEXACT\,
datac => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_RNIFKJL_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011101111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_60_SUM0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_2_C0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(45),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(46),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(14));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(25));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(21),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(117),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datac => \GRLFPC2_0.FPI.LDOP_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011110010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(118),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datac => \GRLFPC2_0.FPI.LDOP_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(50));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(35));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(20));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(40),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(40));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(47));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101000001010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_3\);
\GRLFPC2_0_COMB_V_STATE_1_IV_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010000000")
port map (
combout => \GRLFPC2_0.COMB.V.STATE_1_IV\(1),
dataa => N_19,
datab => \GRLFPC2_0.V.STATE_1_SQMUXA_X\,
datac => CPO_EXCZ,
datad => \GRLFPC2_0.COMB.V.STATE\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_NOTPROP_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100110011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.NOTPROP_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP_1_SUM0_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP_1_C0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_SUM0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_3_RNIDMBD1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110100110010110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN16_NOTPROP_0_S\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_SUM0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_C0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN18_STKGEN_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110100101101001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN18_STKGEN_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP_1_C0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_SUM0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.FPI.LDOP_REP3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(38));
GRLFPC2_0_UN1_FPOP7_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100000")
port map (
combout => \GRLFPC2_0.UN1_FPOP7_1\,
dataa => N_88,
datab => N_87,
datac => \GRLFPC2_0.COMB.FPDECODE.FPOP3_0_A2\,
datad => \GRLFPC2_0.UN1_RS1V_0_SQMUXA_0\);
GRLFPC2_0_COMB_RS1D_1_U: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111011110000000")
port map (
combout => \GRLFPC2_0.COMB.RS1D_1_U\,
dataa => N_76,
datab => \GRLFPC2_0.COMB.RS1_1_SN_M2_I_A2\,
datac => \GRLFPC2_0.COMB.FPDECODE.RS1D5_0_A2\,
datad => \GRLFPC2_0.RS1D_CNST_0_A2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_14: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000111110000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_14\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_11_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_14_A\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_12_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_14_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010101100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_14_A\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_8_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_9_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(19));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_35_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110010001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN14_CONDITIONAL\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_42: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_42\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN18_XZXBUS_37_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_27\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_41: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_41\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN18_XZXBUS_32_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_25\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_38: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_38\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN18_XZXBUS_40_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_19\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_37: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_37\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(35),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN18_XZXBUS_19_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_17\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_36: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_36\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN18_XZXBUS_28_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(45),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_15\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_6\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_11\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_8_0_A2\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_3_1\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1\(26),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_9\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_0_23_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_23\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_16\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_15\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_14\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_17\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_1_19_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_19\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_1\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_0\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_11\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_17\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_23\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_15\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_17\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_16\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_14\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_22\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_0\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_7\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_15\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_19\);
GRLFPC2_0_COMB_WREN125_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.COMB.WREN125_1\,
dataa => \GRLFPC2_0.R.X.LD\,
datab => \GRLFPC2_0.R.I.V\,
datac => \GRLFPC2_0.COMB.ISFPOP2_1_X\,
datad => \GRLFPC2_0.COMB.V.I.EXEC\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN2_NOTDECODEDUNIMP: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110111111101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.STARTSHFT.UN2_NOTDECODEDUNIMP\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(66),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(64),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.STARTSHFT.UN3_NOTDECODEDUNIMP\);
GRLFPC2_0_R_A_RDD_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.R.A.RDD_0_0_G1\,
dataa => \GRLFPC2_0.COMB.RDD_1.M14_0_A2_2_2_X\,
datab => \GRLFPC2_0.COMB.RDD_1.M14_0_A2_3_0\,
datac => \GRLFPC2_0.COMB.RDD_1.M14_0_A2_1_X\,
datad => \GRLFPC2_0.COMB.RDD_1.M14_0_A2_0\);
\GRLFPC2_0_R_STATE_RNO_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100110000000000")
port map (
combout => \GRLFPC2_0.R.STATE_0_0_0__G1\,
dataa => N_19,
datab => \GRLFPC2_0.V.STATE_1_SQMUXA_X\,
datac => CPO_EXCZ,
datad => \GRLFPC2_0.COMB.V.STATE_7_IV_I\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_RNIO4M01: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011101111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_SUM1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_C0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_ADD0\);
GRLFPC2_0_RS1D_CNST_0_A2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.RS1D_CNST_0_A2\,
dataa => N_79,
datab => N_81,
datac => N_88,
datad => \GRLFPC2_0.RS1D_CNST_0_A2_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_OPREXC_RNII87R: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW\(77),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(46),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW_0\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN1_TEMP\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXC\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_6\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_6\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_6\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_7\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_15\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_19\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_16\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_15\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_17\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_9\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_A\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_13\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_12\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_A\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_6\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_8_0\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_11\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_10\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_14\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_12\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_13\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_15\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_7\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_10\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_6\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_12\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_8\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_9\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_7\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_10\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_2\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2_4\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(37),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_1\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_35__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12\(35),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_35__G2_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1_A2\(39),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_35__G2_3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_7\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_9\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_10\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_11\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_15\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_12\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_17\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_16\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_9\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_11\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_21\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_4\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_5_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_9\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_10\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_7\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_12\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_6\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_10\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_3_0_O2\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_2_0_O2\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_4\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_4\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_11\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_10\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_6\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_14\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_7\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_18\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_6\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_7\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_5_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_2_RNIPB7B3_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_8\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_7\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_9\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_11\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_10\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_7\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_5\);
GRLFPC2_0_R_I_V_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110011000100")
port map (
combout => \GRLFPC2_0.R.I.V_1_0_G2\,
dataa => N_17,
datab => \GRLFPC2_0.R.I.V_1_0_G2_0\,
datac => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2\,
datad => \GRLFPC2_0.COMB.UN6_IUEXEC\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTRESETORUNIMP: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111000111110001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.STARTSHFT.UN3_NOTRESETORUNIMP\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(66),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.STARTSHFT.UN3_NOTDECODEDUNIMP\);
GRLFPC2_0_COMB_RS2D_1_IV_0_O2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101000000")
port map (
combout => \GRLFPC2_0.COMB.RS2D_1_IV_0_O2\,
dataa => N_65,
datab => \GRLFPC2_0.COMB.RS2D_1_IV_0_O2_0\,
datac => \GRLFPC2_0.RS1V_0_SQMUXA_1_0_A2_2_X\,
datad => \GRLFPC2_0.COMB.RS2D_1_IV_0_A2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(45),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(45),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(46),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(46),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(16),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(41),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(24),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(25));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(12),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(10),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(21),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(21),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(26),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(14),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(14));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(22),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(23),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(50),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(50));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(39),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(43),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(37),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(35),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(35));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(20),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(20));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(30),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(28),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(15),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(40),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(40),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(40));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_5_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(116),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datac => \GRLFPC2_0.FPI.LDOP_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(0));
GRLFPC2_0_COMB_SEQERR_SEQERR_0_A3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010000000")
port map (
combout => \GRLFPC2_0.COMB.SEQERR.SEQERR_0_A3\,
dataa => \GRLFPC2_0.R.A.SEQERR_RET_3\,
datab => \GRLFPC2_0.RS2_0_SQMUXA_2\,
datac => \GRLFPC2_0.RS2_0_SQMUXA_3\,
datad => \GRLFPC2_0.COMB.SEQERR.UN13_OP\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_233_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111000010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_233__G0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(233),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0\(233),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M2_0\);
GRLFPC2_0_COMB_UN1_V_STATE: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.COMB.UN1_V.STATE\,
dataa => \GRLFPC2_0.COMB.V.STATE_7_IV_I\(0),
datab => \GRLFPC2_0.COMB.V.STATE\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_67_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW_6_0_67__G0_I_O4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.FPI.START\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_71_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110111001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.UN36_PCTRL_NEW_I_0_G0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.UN4_TEMP2\,
datab => \GRLFPC2_0.FPI.START\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.TEMP_25\);
\GRLFPC2_0_R_FSR_FTT_RNO_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010000000")
port map (
combout => \GRLFPC2_0.R.FSR.FTT_0_0_0__G1\,
dataa => N_8,
datab => \GRLFPC2_0.R.FSR.FTT\(0),
datac => \GRLFPC2_0.UN1_FPCI_21\,
datad => \GRLFPC2_0.N_1570_I_I_A2\);
\GRLFPC2_0_R_FSR_FTT_RNO_0_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101110111011")
port map (
combout => \GRLFPC2_0.R.FSR.FTT_0_0_2__G1_A\,
dataa => \GRLFPC2_0.COMB.UN1_FPCI_X\,
datab => \GRLFPC2_0.R.X.SEQERR\,
datac => \GRLFPC2_0.R.FSR.FTT\(2),
datad => \GRLFPC2_0.UN1_FPCI_21\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(38));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_234_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111000010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_234__G0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(234),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0\(234),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_232_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111000010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_232__G0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(232),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0\(232),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M2_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_16_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G_32\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD12\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.REEXCOVUV.UN20_LOCOV\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_4510_A2_7\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_18_2\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1_A2_0\(39),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2\(38));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_51_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN14_CONDITIONAL\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIKT3S_315_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111100101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(315),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1_1_A\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNINI7K_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110100000000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1_1_A\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN6_NOTPROP_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_33: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010000101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_33\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(47),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(47));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_32: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001001001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_32\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(53));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_31: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010000101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_31\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(56));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_30: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010000101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_30\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(21),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(36));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_29: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010000101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_29\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(38),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(22),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(22),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(38));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_27: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010000101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_27\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(46),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(20),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(20),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(46));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_25: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001001001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_25\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(42));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_24: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010000101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_24\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(26),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(51));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_23: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010000101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_23\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(43),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(43));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_22: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001001001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_22\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(49),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(41));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_21: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001001001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_21\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(24),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(24));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_19: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001001001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_19\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(54));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_17: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010000101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_17\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(39),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(23),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(39));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_15: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010000101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_15\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(44));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_12: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001001001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_12\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(15),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(14));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001001001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_6\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010000101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZZERO_1_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(12),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110110110111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_9\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110110110111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_5\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(8));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111000010110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_2_RNIDEGV_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_10\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_2\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_3_0_O2\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_9\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_0_0_O2\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_22\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_12\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_13\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_18\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_20\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_15\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_24\(58),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_7\(58),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_14\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_12\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_4\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_2\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_7\(62),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_9\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_1_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_0_I_O2\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_9_0_A2\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_0_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_16\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_6\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_12\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_7\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_14\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_4\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_0\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_7\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_11\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_11\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_0_A2\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_0_A2_0\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_7\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_21_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_21\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_11\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_11\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_16\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_10\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_20_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_20\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A2_9\(47),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_9_TZ\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_7\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_14\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_1_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_12\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A19\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_1\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_3_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_14\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_5\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_17\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12\(20),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_10\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_17\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_18\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_1\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_7\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_13\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_18\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_4\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_11\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_15\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_1_17_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_17\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_3_TZ\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_15_2\(60),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_3_0\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_13\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_23\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_18\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_1\(60),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_8\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_19\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_0_RNIJJGV6_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_24\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_11_0_A2\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_20\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_15\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_24_RNI9COG1_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_23\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_24\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_7\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_11\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_18\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_20\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_11\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_9\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_8\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_10\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_19\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_9\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_16\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_15\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_19\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_6\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_11\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_17\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_21\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_3\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_14\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_18\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_17\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_21\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_20\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_6\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_13\);
GRLFPC2_0_UN1_RS1V_0_SQMUXA_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100100000")
port map (
combout => \GRLFPC2_0.UN1_RS1V_0_SQMUXA_0\,
dataa => N_68,
datab => N_63,
datac => \GRLFPC2_0.RS1V_0_SQMUXA_1_0_A2_0_3\,
datad => \GRLFPC2_0.RS1V_0_SQMUXA_1_0_A2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTDECODEDUNIMP: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.STARTSHFT.UN3_NOTDECODEDUNIMP\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(67),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.ENTRYPOINT_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.STARTSHFT.UN3_NOTDECODEDUNIMP_A\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTDECODEDUNIMP_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100011111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.STARTSHFT.UN3_NOTDECODEDUNIMP_A\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_1_1\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN1_S\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.ENTRYPOINT_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_GRFPUF_0_RNIDSD8_0_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110011111000011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_374__G0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF_0\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF_0\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_374__G0_A\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_2_RNIQRG7_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000101000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_374__G0_A\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF_0\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF_0\(0));
GRLFPC2_0_R_A_LD_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC2_0.R.A.LD_0_0_G1\,
dataa => \GRLFPC2_0.R.A.LD_0_0_G1_2_X\,
datab => \GRLFPC2_0.R.A.LD_0_0_G1_3\,
datac => CPO_EXCZ,
datad => \GRLFPC2_0.N_939_I_I_A2\);
GRLFPC2_0_FPI_START: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC2_0.FPI.START\,
dataa => N_17,
datab => \GRLFPC2_0.R.MK.RST2\,
datac => \GRLFPC2_0.COMB.V.MK.RST_1_0_A2\,
datad => \GRLFPC2_0.R.A.FPOP_0_0_G1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN11_WQSTSETS\);
GRLFPC2_0_V_STATE_2_SQMUXA_I_A2_0_RNIJV401: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010110000")
port map (
combout => \GRLFPC2_0.COMB.V.STATE\,
dataa => \GRLFPC2_0.COMB.UN1_FPCI_X\,
datab => \GRLFPC2_0.R.X.SEQERR\,
datac => \GRLFPC2_0.COMB.V.STATE_0\,
datad => \GRLFPC2_0.V.STATE_2_SQMUXA_I_A2_0\);
GRLFPC2_0_COMB_V_I_EXEC_4_IV_0_A2_X_RNIDL351: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010101000")
port map (
combout => \GRLFPC2_0.N_1570_I_I_A2\,
dataa => \GRLFPC2_0.R.I.V\,
datab => \GRLFPC2_0.COMB.V.I.EXEC_4_IV_0_A2_X\,
datac => \GRLFPC2_0.R.I.RDD_0_0_G1_0_8238_I_O4\,
datad => \GRLFPC2_0.COMB.UN1_MEXC_1\);
GRLFPC2_0_COMB_UN3_IUEXEC_RNI9GFG3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.N_939_I_I_A2\,
dataa => N_89,
datab => N_90,
datac => \GRLFPC2_0.N_939_I_I_A2_0_1_X\,
datad => \GRLFPC2_0.N_939_I_I_O2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_3_1\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_11_0_A2\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_10_1\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_0\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O6_3_RNIARA81_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_30__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_2\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O6_3\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_30__G2_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_30__G2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A7\(29),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_0\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_14\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_7\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_24__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2\(24),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_1\(24),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(24),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_23__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_23__G2_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_23__G2_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_22__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_0_I_O2\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_1_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2\(22),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_15__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(38),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_4_0_A2\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_15__G2_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_15__G2_3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_RNI6U5H_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_8__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_1_0_A2\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_18_2\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A7_0\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O7_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_1__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN1_S_DYADIC_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_0_A2\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1\(1));
GRLFPC2_0_R_X_SEQERR_RNI5TGU1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001000")
port map (
combout => \GRLFPC2_0.R.I.V_1_0_G2_0\,
dataa => \GRLFPC2_0.R.I.V_1_0_G2_0_0_X\,
datab => \GRLFPC2_0.R.I.V_1_0_G2_0_3\,
datac => \GRLFPC2_0.ANNULRES_0_SQMUXA_10\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_XX_RNIT1JJ_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001111110010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_YY_RNIVK6I_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100100001001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_6_M3_E\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_YY\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_XX_RNISTIJ_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001111110010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_YY_RNIJK6I_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100100001001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_4_M3_E\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_YY\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_3_M4_I_X2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100011000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_3_M4_I_X2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_3_M1_E_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_3_M4_I_X2_A\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_3_M4_I_X2_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_3_M4_I_X2_A\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI05LB_0_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP_1_C0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(370),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_1_RNII4B9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_2_C0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI85LB_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_C0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(369),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.CIN_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIU51B_0_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_C0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.TEMP2_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN18_XZXBUS_13_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001100110011001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN18_XZXBUS_13_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111010111100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111010111100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111010111100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111010111100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111010111100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111001010100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111001010100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111010111100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_GRFPUF_0_RNIDSD8_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_375__G0_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF_0\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF_0\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_374__G0_A\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111010111100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(9));
\GRLFPC2_0_COMB_V_STATE_7_IV_I_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110100")
port map (
combout => \GRLFPC2_0.COMB.V.STATE_7_IV_I\(0),
dataa => \GRLFPC2_0.COMB.UN1_FPCI_X\,
datab => \GRLFPC2_0.R.X.SEQERR\,
datac => \GRLFPC2_0.R.STATE\(0),
datad => \GRLFPC2_0.V.STATE_2_SQMUXA_I_A2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_A\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_A_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010000000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_A\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(43),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M14\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110110001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19_3_0_.M4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_SN_M3_E\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_SN_M3_E\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19_3_0_.M3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_SN_M3_E\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19_3_0_.M2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_12_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_12_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN14_CONDITIONAL\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_OPREXC: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111101111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXC\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN14_CONDITIONAL\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2\(37),
dataa => N_34381_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_18_2\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2\(38));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOINSTANDNOEXC_1_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001100100011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.UN4_TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.TEMP_25\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110110110111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(12),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_10_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000111110011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN5_SHDVAR\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN19_GEN_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111100001111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_SUM1_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_SUM0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_2_0_O2_RNIL4U31_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_8\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_0_A2\(41),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_1_2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_2_0_O2\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_3_RNIG3BB_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_6\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_11_0_A2\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_3\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_2\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_4_0_A2\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_18\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\(58),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O29_6\(58),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_11\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_17\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_1\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_11\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_10\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_16\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_3\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_1\(58),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_11\(58),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_4\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_14\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A22_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_26_2\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_0\(58),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_10\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_10\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_30\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_16_1\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_4\(50),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_13\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_4\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_3\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_16\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_8\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_12\,
dataa => N_33157_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_14_0\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_6\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_14\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7_2\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_12_0_A2\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_12\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_8\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_7\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_16\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_11\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_13\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_10\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_15\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_5\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_12\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_O2\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_9_0_A2\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(28),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_11\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_5_0\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_3\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_9\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_13\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_2\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_1\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_8\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_10\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_11_0_A2\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_10_1\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_0\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_6\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_11\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_3_I_O2\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_9_0_A2\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_10\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_3\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_1\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_9\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A18\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_16\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_14_0_A2\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_5\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_8\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_5\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_3_TZ\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_7\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_6\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_19_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_19\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_14_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_4\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_4\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_19_A\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_19_A_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_19_A\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A7_1\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_9_1\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_20_2\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_14\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_18_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_18\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN1_S_DYADIC_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_1_TZ\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_0\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_12\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_19\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_16\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_9\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_12\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100011111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_18\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_6_1\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_3_1\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_18_A\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_18_A\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(13),
datab => N_28871_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_26\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_5_2\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_17\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_22\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_1\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_6\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_15\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_3_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_10\,
dataa => N_34483_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_16_1\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_2\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_4\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_12\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_4\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_5\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A20\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_6\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_10\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_4_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O20_5\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_4\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_9\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_7\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_13\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_3\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_12\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_15\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_1_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_13\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_2_2\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_17_1\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_13\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_6\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_0_18_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_18\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80),
datab => N_33157_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_M2_0\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_12\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_0_17_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_17\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_11\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_17_2\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_11\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_10\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_0_16_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_16\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_23_0\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_7_2\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_0\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_0\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_0_15_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_15\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_25_0\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_25_1\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_A28\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_7\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_10\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A15_0\(18),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_5\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_2\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_7\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_9\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_1\(18),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_14_0_A2\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_2_RNICPPA_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_8\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_5\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_6\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_10_0_RNIMJUP_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_10_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_14_0_A2\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_15\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_0_A2\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_14\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A22_0\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_6\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_5\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_8\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_1_14_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_14\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_1\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_7\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_6\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_1_13_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_13\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_1_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_5\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_8_1\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_4\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_O2\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_9_0_A2\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_0_A2\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_0_A2_0\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_22\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_5\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_2\(60),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_22\(60),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_17\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_21\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O25\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_3_1\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_15\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_20\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1_A2_1_1\(39),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_26_2\(60),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_12\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_11_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_19\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_12\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30\(60),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_3\(60),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_10\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_6\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_2_2\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_2_3\(62),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_21_RNIHLDS5_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_20\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_0\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_21\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_1\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_13\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_2_RNI078L_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_18\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_12\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_2\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_9\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_3\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_15\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_14_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_1_2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_11\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_7\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_17\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_17\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_19\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_12\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_15\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O21_3\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7_0\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_5\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_9\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_19\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_6_2\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_6_1\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_0\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_12\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_18\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_3\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_16\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_6\(60),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_16\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A27\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_2\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_23\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_9\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_9_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_18\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_22\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_7\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_12\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_16\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_I_A26_1\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_16\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_16_A\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100111100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_16_A\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_10_1\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_2\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_19\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_11\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_8\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_13\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_18\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_5\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_6\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_8_0_A2\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_11_0_A2\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_4\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_10\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_8_1\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_2_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_13\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_6\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_15\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_1\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_10_2\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_10\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_14\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_7\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_1\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A21\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_13\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_13\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_15_3\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_15_4\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_6\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_7\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_12\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_18\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_9\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_16\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_16\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_4\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_12\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_15\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_22\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_28\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_10\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101000110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_8\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_0_2\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_0_I_O2\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_9_0_A2\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_5_TZ\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_0\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_1_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_8732\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_10\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O16\(49),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_1_1\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_0_A2_0\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_5\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_9\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_6\(49),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_10\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_11\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_2\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_8\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_1_1\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_9_1\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A16\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_1_1\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_8_1\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_16_1\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_16_4\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_8715\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A13\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_5\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_12_0\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_12_0_0\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_14\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_0\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_1_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_1_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_5_1\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_0_1\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_0_A2_0\(28),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_0_A2\(28));
GRLFPC2_0_R_I_EXEC_RNI62DN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111111011100")
port map (
combout => \GRLFPC2_0.R.I.V_1_0_G2_0_3\,
dataa => \GRLFPC2_0.COMB.UN1_FPCI_X\,
datab => \GRLFPC2_0.R.I.EXEC\,
datac => \GRLFPC2_0.R.X.FPOP\,
datad => \GRLFPC2_0.R.I.V_1_0_G2_0_3_A\);
GRLFPC2_0_COMB_UN1_FPCI_1_X_RNIP4V8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101011111")
port map (
combout => \GRLFPC2_0.R.I.V_1_0_G2_0_3_A\,
dataa => \GRLFPC2_0.COMB.UN1_FPCI_1_X\,
datab => \GRLFPC2_0.COMB.UN1_FPCI_2_X\,
datac => \GRLFPC2_0.R.M.FPOP\,
datad => \GRLFPC2_0.R.E.FPOP\);
GRLFPC2_0_COMB_WREN1_9_IV_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC2_0.COMB.WREN1_9_IV_0\,
dataa => \GRLFPC2_0.COMB.WREN1_9_IV_0_A\,
datab => \GRLFPC2_0.R.X.SEQERR\,
datac => \GRLFPC2_0.R.X.LD\,
datad => \GRLFPC2_0.R.X.AFSR\);
GRLFPC2_0_COMB_WREN1_9_IV_0_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010110001")
port map (
combout => \GRLFPC2_0.COMB.WREN1_9_IV_0_A\,
dataa => N_353,
datab => N_358,
datac => \GRLFPC2_0.COMB.WREN12_X\,
datad => \GRLFPC2_0.COMB.UN1_FPCI_X\);
GRLFPC2_0_RS1D_CNST_0_A2_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010100010100000")
port map (
combout => \GRLFPC2_0.RS1D_CNST_0_A2_0\,
dataa => N_78,
datab => \GRLFPC2_0.RS1D_CNST_0_A3_0_A2_1_X\,
datac => \GRLFPC2_0.RS1D_CNST_0_A3_0\,
datad => \GRLFPC2_0.RS1D_CNST_0_A3_0_A2_0_0\);
GRLFPC2_0_COMB_WREN2_9_IV_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC2_0.COMB.WREN2_9_IV_0\,
dataa => \GRLFPC2_0.COMB.WREN2_9_IV_0_A\,
datab => \GRLFPC2_0.R.X.SEQERR\,
datac => \GRLFPC2_0.R.X.LD\,
datad => \GRLFPC2_0.R.X.AFSR\);
GRLFPC2_0_COMB_WREN2_9_IV_0_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001001110")
port map (
combout => \GRLFPC2_0.COMB.WREN2_9_IV_0_A\,
dataa => N_353,
datab => N_358,
datac => \GRLFPC2_0.COMB.WREN12_X\,
datad => \GRLFPC2_0.COMB.UN1_FPCI_X\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_14\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_15\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.NOTAM2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_27\);
GRLFPC2_0_COMB_RS2D_1_IV_0_A2_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC2_0.COMB.RS2D_1_IV_0_A2_0\,
dataa => N_66,
datab => N_76,
datac => N_69,
datad => \GRLFPC2_0.COMB.RDD_1.M14_0_O2\);
GRLFPC2_0_COMB_PEXC8_RNI47GK2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC2_0.R.A.FPOP_0_0_G1\,
dataa => \GRLFPC2_0.COMB.RS1_1_SN_M2_I_A2\,
datab => \GRLFPC2_0.N_939_I_I_2_X\,
datac => CPO_EXCZ,
datad => \GRLFPC2_0.COMB.FPOP_0_0_O2\);
GRLFPC2_0_COMB_RDD_1_M14_0_A2_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.COMB.RDD_1.M14_0_A2_0\,
dataa => \GRLFPC2_0.COMB.RS1_1_SN_M2_I_A2\,
datab => \GRLFPC2_0.COMB.RDD_1.M14_0_O2\,
datac => \GRLFPC2_0.COMB.FPDECODE.RS1D5_0_A2_0\,
datad => \GRLFPC2_0.RS1V_0_SQMUXA_1_0_A2_1_X\);
GRLFPC2_0_COMB_UN6_IUEXEC: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.COMB.UN6_IUEXEC\,
dataa => \GRLFPC2_0.R.MK.RST2\,
datab => \GRLFPC2_0.COMB.UN3_IUEXEC\,
datac => \GRLFPC2_0.COMB.V.MK.RST_1_0_A2\,
datad => \GRLFPC2_0.COMB.UN6_IUEXEC_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPBREGLOADEN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datac => \GRLFPC2_0.FPI.LDOP_REP0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLAREGEXP.EXPAREGLOADEN_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_3_0_O2_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_3_0_O2\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7_2\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_12_0_A2\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_26\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_27\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1_A2_1_1\(39),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_1_0_A2\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_4\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1_A2\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_1_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100011111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_1\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_0_A2\(41),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_3_1\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_1_0\(38));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_14\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_4_0_A2\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_2\(22),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(22),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_1\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_44__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_18_2\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_1_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_44__G2_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_12_I_O2_RNILM641_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110111111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_12_I_O2\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_14\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100011111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_14__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_4785_A2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_9_0_A2\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_14__G2_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_2__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_1_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_45\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_9__G2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_XX_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000011011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN25_NOTXZYFROMD\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_7_M3_E_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_XX_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000011011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN25_NOTXZYFROMD\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_5_M3_E_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP2\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN14_CONDITIONAL: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN14_CONDITIONAL\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_4\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_5\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN3_NOTAZERODENORM\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001000011101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_13_M1_E\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.EXTEND.TEMP_1\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN18_XZXBUS_18_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001100110011001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN18_XZXBUS_18_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(18),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(18));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN18_XZXBUS_28_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001100110011001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN18_XZXBUS_28_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(28));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN18_XZXBUS_37_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011110000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN18_XZXBUS_37_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14_171_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_14\(171),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_T_3\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN18_XZXBUS_19_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001100110011001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN18_XZXBUS_19_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(45),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP2\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(45),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(46),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP2\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(46),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP2\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010010111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(16),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(35));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000011111011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP2\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(39),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8_A\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_A_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100001111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8_A\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(40),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010010111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(16),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010010111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(23),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(12),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000011111011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8_A\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_A_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100001111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8_A\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000011111011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(24),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8_A\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_A_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100001111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8_A\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010010111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(10),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(14),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010010111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(20));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(21),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(21),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(20));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(22),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(23),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP2\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(50),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP2\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(50));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP2\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP2\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP2\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP2\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP2\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000011111011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP2\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(40),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8_A\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_A_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011110001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8_A\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP2\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(43),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010010111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP2\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000011111011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP2\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(37),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8_A\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_A_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100001111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8_A\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP2\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(35),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(15),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(14));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000011111011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(40),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP2\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8_A\(40));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_A_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011110001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8_A\(40),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(40),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000011111011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8_A\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_A_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011110001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8_A\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000011111011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(26),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8_A\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_A_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011110001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8_A\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(28),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000011111011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8_A\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_A_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100001111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8_A\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(28),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111001010100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP2\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP2\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN2_DIVMULTV_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_DIVMULTV\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF_0\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF_0\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF_0\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF_0\(0));
GRLFPC2_0_COMB_UN3_IUEXEC_RNI61LG2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111010100000")
port map (
combout => \GRLFPC2_0.N_939_I_I_O2\,
dataa => \GRLFPC2_0.N_939_I_I_A2_1_0\,
datab => \GRLFPC2_0.N_939_I_I_A2_0_0\,
datac => \GRLFPC2_0.COMB.FPOP_0_0_O2_0_2\,
datad => \GRLFPC2_0.COMB.UN3_IUEXEC\);
GRLFPC2_0_COMB_SEQERR_UN13_OP: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.COMB.SEQERR.UN13_OP\,
dataa => \GRLFPC2_0.R.A.AFQ_RET\(7),
datab => \GRLFPC2_0.R.A.MOV_RET\(15),
datac => \GRLFPC2_0.COMB.SEQERR.UN13_OP_A\,
datad => \GRLFPC2_0.N_782\);
GRLFPC2_0_COMB_SEQERR_UN13_OP_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001100000001")
port map (
combout => \GRLFPC2_0.COMB.SEQERR.UN13_OP_A\,
dataa => \GRLFPC2_0.R.A.MOV_RET\(12),
datab => \GRLFPC2_0.R.A.MOV_RET\(13),
datac => \GRLFPC2_0.R.A.AFQ_RET\(5),
datad => \GRLFPC2_0.R.A.MOV_RET\(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPAREGLOADEN\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datac => \GRLFPC2_0.FPI.LDOP_REP0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLAREGEXP.EXPAREGLOADEN_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_233_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0\(233),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233),
datac => \GRLFPC2_0.FPI.LDOP_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLAREGEXP.EXPAREGLOADEN_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN18_XZXBUS_40_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011110000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN18_XZXBUS_40_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(40));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN18_XZXBUS_32_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011110000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN18_XZXBUS_32_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN2_MIXOIN_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111100001101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(371),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_A\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN2_MIXOIN_A_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001011100010111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_A\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_RNIIE0U_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000111101110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN10_NOTPROP_0_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP_1_SUM0_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000011111011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8_A\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_A_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100001111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8_A\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(10));
GRLFPC2_0_R_I_RDD_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011001010")
port map (
combout => \GRLFPC2_0.R.I.RDD_0_0_G1_0_8238_I\,
dataa => \GRLFPC2_0.R.I.RDD\,
datab => \GRLFPC2_0.R.X.RDD\,
datac => \GRLFPC2_0.R.I.RDD_0_0_G1_0_8238_I_O4\,
datad => \GRLFPC2_0.R.I.RDD_0_0_G1_0_8238_I_A3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_8\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP2\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(37));
GRLFPC2_0_COMB_V_I_EXEC_4_IV_0_A2_X_RNIQ3AU1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111000001110")
port map (
combout => \GRLFPC2_0.COMB.V.I.EXEC\,
dataa => \GRLFPC2_0.COMB.V.I.EXEC_4_IV_0_A2_X\,
datab => \GRLFPC2_0.R.I.RDD_0_0_G1_0_8238_I_O4\,
datac => \GRLFPC2_0.N_1570_I_I_A2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_232_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0\(232),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(232),
datac => \GRLFPC2_0.FPI.LDOP_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLAREGEXP.EXPAREGLOADEN_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_234_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000010101010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0\(234),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.FPI.OP2_X\(62),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPAREGLOADEN_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN20_LOCOV: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101110111011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.REEXCOVUV.UN20_LOCOV\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD11\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN30_CONDITIONAL_M5\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_0_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_0\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_1\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_7\(38),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_4\(37));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100110011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(4));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_2_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_3_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_17_0_A2_RNI7GIG_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100011111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_16__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_1_0\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_A26_17_0_A2\(60),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0_0\(10),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_0\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110010100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_2_0\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_11\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_9_0_A2\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_23\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_5\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_2_2\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_5_1\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_34_2\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_1_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_4_0\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_2_0_I_O2\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_1_0_A2\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_5\(25));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_17_2\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_0\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_4\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_13\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_1_1\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_9023_TZ\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_6\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_5\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_12\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_21\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_25\(58),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_6\(58),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_23\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_12_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_11\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_2\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_1\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_2_1\(58),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_10\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_19_0\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A25_1\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_18\(58),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_9\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_4_1\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_12_0_A2\(62),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_6\(50));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_A2_1\(26),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000011111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_6\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_7_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_2_0_A2\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_6_A\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_6_A\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0_2\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_2_0\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_2_0_I_O2\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_14\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101011000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_6_1\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_25_1\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_1_0\(50),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_3_1\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_11\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_8\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_10_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O21\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_7\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_10\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_17_1\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A13_1\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_16_4\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_0\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_9\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_5_0\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_26_2\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_20\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_8\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_18\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_6\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_2\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_10\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_6\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0_1\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_9_3\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_8\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_0_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_A28_11_0_A2\(47),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_9_7495\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_8_1\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_2_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_0_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_11_0_A2\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_14_2\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_2_0_A2\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_1\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_10\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O21_2\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_1_1\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A21\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_2\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_3_1\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_8\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_1_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_0_2\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_14\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_12_2\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_2_0_A2\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_2\(44),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_6\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_6\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_1_0_A2\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11_2\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_4\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_5\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_25\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_17_1\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_4_2\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_4785_A2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_14_2\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_1\(7),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_16_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_16\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A22_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_M27\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_8_2\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_14_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_14\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_3_0\(47),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_1\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_14_A\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_14_A_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_14_A\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN1_S_DYADIC_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_I_A26_1\(31),
datac => N_29496_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_7\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_12_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_12\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_5_0\(47),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_X2_0\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_2\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_0\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_10_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_10\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A2_9\(47),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_9_7495\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_6_1\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_16\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_7_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_7\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_16_1\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_6\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_9_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_16\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_2_2\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_2_0\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A28\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_11\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_11_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_14\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_0_0\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_10\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_4\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_12\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_10_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_5\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_8\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_3\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_0_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_10\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_6\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_8\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_5\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_2_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_6\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A19_2\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_1\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_6\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_8\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_1\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_6\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_19\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_10_1\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_2\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_12\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11_0\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11_2\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_5\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_11\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7_0\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7_2\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_2\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110010100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_9_0\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_8\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_4_2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_0_1\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_9_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_6\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A28_1\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_4_1\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_11\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_0_14_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_14\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_2\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_18_3\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_16\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_6\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_0_13_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_13\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_22\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_15\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_17\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_24\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_0_12_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_12\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_O28_6\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_10_1\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_19\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_14\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_0_10_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_10\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A28_1\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_4_2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_11_0\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_1\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_3_0\(18),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_3_1\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_6\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_0\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_20_2\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_4\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_2\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_11\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_11_0\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_9\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_0_A2_0\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_1_11_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_11\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_2\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_O24_3\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_5_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_2\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000011111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_1_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2_3_A\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001101011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2_3_A\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_17_2\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_2_0_A2\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_12_0_A2\(62),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_26_2\(60));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_0\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_0_I_O2\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000011111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_17\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_5_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_17_A\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_12_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011111100010101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_17_A\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_8692_TZ\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A22_1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_15_2\(60),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O13_0\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_9_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_15\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_21_0\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_7\(60),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_6\(60));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_12\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_4_2\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_16\(60),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_13\(60));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_5\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_2_TZ\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_1\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_0_1\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_0_0\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_6\(62),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_13\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_12_0_RNI958Q_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_17\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_12_0\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_15_4\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_8\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_7\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_20_4_RNITLEL_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_16\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A13_1\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_20_4\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_4\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_6\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_X2_RNITRLP_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_15\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_3_1\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_6_0\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_4\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_10_1_RNI8MVA5_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100111000001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_13\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_16_1\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_10_1\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_13_A\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_2_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_4_2_RNILUF15_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111001101111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_13_A\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_4_2\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_16_RNIAASF_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_11\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_14_3\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_6_1\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_16\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_5\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_13\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1_A2_1_1\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_12\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O18_4\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_1_1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_17\(60),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_11_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_10\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A19_1\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_13_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_9_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_9\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_9_1\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_7_1_0\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_13_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A25\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_10_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_8\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_14_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_3_0\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_6\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_19\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_12_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_1_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_10_1\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O25\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_2\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_5\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_18_1\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_1\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_1\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_10_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_12\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_9\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_19\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_16\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_3\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_11\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_6\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O18_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_9\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_7_1\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O23\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_13_0\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_0\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_5\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_13_1\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_2_2\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_1\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_17\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_15\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_19\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_24\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_11\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_15\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_17_1\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_2\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_8\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_14\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O27_10\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A28_1\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A3_3_2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_12\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_15_0\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_5\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_5\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_15__G2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_4785_A2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_1_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_11_0_A2\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_0_A2\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101011000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_5_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_25\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_5_TZ\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_A2_1\(26),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_5_0_A2\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_14_2\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_0_I_O2\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_9\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_12\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11_2\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_1\(26),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_14\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_23\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_9\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_8\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_0\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_11_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_12\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_16_1\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_2_TZ\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_18\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_5\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111101010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_11\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_10\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_4_0\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_14_1\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_15\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_18_3\(47),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_23_0\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_17\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_8\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_11_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_13\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_16_0\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_12\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_10\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80),
datab => N_33495_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_2_1\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A26\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_9\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X3\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_24_3\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_3\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_10_1\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\(58),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_1\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101010111000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_12\(60),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_2\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_13\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_6_I_O2\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_2_0_A2\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_7\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_9\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_12_2\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O2\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_4\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_4\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_8\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_1\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O17_1\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_1_2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A17_1\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_2\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_7_A\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_5\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_7_A\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_2\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_20\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000011111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_6\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN1_S_DYADIC_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_6_A\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011110111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_6_A\,
dataa => N_28709_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_3_1_0\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_10\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_18\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_1_1\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_17_0\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_7\,
dataa => N_34483_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0_1_0\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_3\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_14\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_9_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_13\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_34_2\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_18\(60),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_7\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_12\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_5\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A22_1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_26_2\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_29\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_10\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_11\(53),
datac => N_29496_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_6\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_24_1\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A26_1\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_36\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_35__G2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_18_1\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_2_3\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1_A2_1\(39),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_2\(35));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_35__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11_2\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\(58),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1_A2_0\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_6\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_12\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_9\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_4\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_5_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_11_0\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_11_1_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_10\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_5\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datab => N_28871_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_4_1\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_13\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_20_0\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_2_1\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_15\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000101011111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_23__G2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_12\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_23__G2_2_A\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000111110011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_23__G2_2_A\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_10_1\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_3_1\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_O2\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_14\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111001101010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_23__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_O28_5\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_0_I_O2\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_30\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_1_0\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_1_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_1\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_O2\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_1\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A6_3_RNID0LC_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_30__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_3_1\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O6_2\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O25\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A6_3\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A6_2_RNI6TEH_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_30__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A13_1\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O6_1\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_8_1\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A6_2\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_4_0\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_2\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_3\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_0\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X3\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_2_4\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_1_1\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O7_1\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O25\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_3\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_9_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O7_0\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_4\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_1_0_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_1_0\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_37\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_0_2\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_25_1\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_30\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_0_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_14__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_14_2\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11_2\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2\(14),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2\(2));
GRLFPC2_0_R_X_AFQ_RNI44GM: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111100000000")
port map (
combout => \GRLFPC2_0.COMB.V.STATE_0\,
dataa => \GRLFPC2_0.COMB.UN1_FPCI_X\,
datab => \GRLFPC2_0.R.STATE\(0),
datac => \GRLFPC2_0.R.X.AFQ\,
datad => \GRLFPC2_0.R.STATE\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_27: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_27\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_16\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_17\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_24\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_23\);
GRLFPC2_0_RS1V_0_SQMUXA_1_0_A2_0_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.RS1V_0_SQMUXA_1_0_A2_0_3\,
dataa => N_62,
datab => \GRLFPC2_0.COMB.FPDECODE.ST_0_A2_0_A2_0_X\,
datac => \GRLFPC2_0.COMB.FPDECODE.FPOP3_0_A2_1_X\,
datad => \GRLFPC2_0.RS1V_0_SQMUXA_1_0_A2_0_1\);
GRLFPC2_0_COMB_RDD_1_M14_0_A2_3_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.COMB.RDD_1.M14_0_A2_3_0\,
dataa => N_63,
datab => \GRLFPC2_0.COMB.RS1_1_SN_M2_I_A2\,
datac => \GRLFPC2_0.COMB.RDD_1.M14_0_O2_0_X\,
datad => \GRLFPC2_0.COMB.RDD_1.M14_0_A2_2_1\);
GRLFPC2_0_FPI_LDOP: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.FPI.LDOP\,
dataa => \GRLFPC2_0.RIN.MK.LDOP_7\,
datab => \GRLFPC2_0.RIN.MK.LDOP_8\,
datac => \GRLFPC2_0.RIN.MK.LDOP_9\,
datad => \GRLFPC2_0.FPI.LDOP_0_X\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI85LB_0_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010110111010010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_57_SUM0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(369),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.CIN_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIU51B_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001010101101010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_56_SUM0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.TEMP2_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(5));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN26_NOTAINFNAN_4_RNIC5AQ: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111011100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN26_NOTAINFNAN_4\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN26_NOTAINFNAN_5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN4_NOTAINFNAN\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI05LB_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010110111010010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP_1_SUM0_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(370),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_1\);
GRLFPC2_0_R_I_RDD_RNO_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.R.I.RDD_0_0_G1_0_8238_I_A3\,
dataa => \GRLFPC2_0.R.E.FPOP_0_0_G1_X\,
datab => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_13_3\,
datac => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_13_4\,
datad => \GRLFPC2_0.R.I.RDD_0_0_G1_0_8238_I_A3_1\);
GRLFPC2_0_COMB_UN2_HOLDN_0_A2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2\,
dataa => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_0_X\,
datab => \GRLFPC2_0.RS2_0_SQMUXA_3\,
datac => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_11\,
datad => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_13\);
\GRLFPC2_0_R_I_EXC_RNO_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001000")
port map (
combout => \GRLFPC2_0.R.I.EXC_2_0_4__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(41),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.EXCEP_1_TZ\(4),
datac => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN11_WQSTSETS: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000110010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN11_WQSTSETS\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD5\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN4_NOTSHIFTCOUNT1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN9_WQSTSETS_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\);
GRLFPC2_0_COMB_ANNULFPU_1_U_0_O2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110100")
port map (
combout => \GRLFPC2_0.COMB.ANNULFPU_1_U_0_O2\,
dataa => \GRLFPC2_0.COMB.UN1_FPCI_X\,
datab => \GRLFPC2_0.R.X.SEQERR\,
datac => \GRLFPC2_0.COMB.ANNULFPU_1_U_0_O2_1\,
datad => \GRLFPC2_0.COMB.ANNULFPU_1_U_0_O2_0\);
GRLFPC2_0_V_STATE_2_SQMUXA_I_A2_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011001000")
port map (
combout => \GRLFPC2_0.V.STATE_2_SQMUXA_I_A2_0\,
dataa => \GRLFPC2_0.R.I.EXEC\,
datab => \GRLFPC2_0.R.I.V\,
datac => \GRLFPC2_0.R.I.RDD_0_0_G1_0_8238_I_O4\,
datad => \GRLFPC2_0.COMB.UN1_MEXC_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN26_NOTBINFNAN_RNIBOPJ: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000010101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN3_NOTBZERODENORM\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN26_NOTBINFNAN\);
GRLFPC2_0_RS1V_0_SQMUXA_1_0_A2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.RS1V_0_SQMUXA_1_0_A2\,
dataa => \GRLFPC2_0.COMB.FPDECODE.ST_0_A2_0_A2_0_X\,
datab => \GRLFPC2_0.COMB.FPDECODE.FPOP3_0_A2_1_X\,
datac => \GRLFPC2_0.RS1V_0_SQMUXA_1_0_A2_3_X\,
datad => \GRLFPC2_0.RS1V_0_SQMUXA_1_0_A2_2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_RNO_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_115__G0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_115__G0_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(115),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(115),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN10_U_SNNOTDB_1_RNIJK0S: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100111110101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.UN10_U_SNNOTDB_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.TOGGLESIG\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_2_0_O2_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_2_0_O2\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_A2_1\(26),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_2_0_O2_0\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A28_4_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_4\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A22_1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_M2\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A13_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_10\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_47__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_25_1\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_22\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_9\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_14\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_41__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_37\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_1_0_A2\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2\(40),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(38));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000011111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_21__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_4_1\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_1_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_21__G2_A\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010100111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_21__G2_A\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_22_1\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_2_0_A2\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_26_2\(60),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_5_0_A2\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_11_RNIM9ER_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_1\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_11\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_4_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_0_2\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_4_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_3_TZ_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_RNIJBEG_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100100111001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(12),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_RNIHBEG_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100100111001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_YY_RNIJJOK_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100100001001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_YY\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_YY_RNIAAJJ_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100100001001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_YY\(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_114_RNI68NL: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010010111000011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_95_RNI6DFD: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110000011110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM_A\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_8732\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_0_0\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_7_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010100010100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_8715\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_O13\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_18_1_0\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_17_1\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_20__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7_2\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11_2\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_3_1\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12\(20));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.EXTEND.TEMP_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_1_RNII4B9_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001010101101010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_2_SUM0_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_SA_I_1_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001010101101010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.SA_I_1_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.TEMP2_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001000011101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(14),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(14),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001000011101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(15),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001000011101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(16),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010000011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010000011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010000011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(20),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(20),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010000011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(23),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010000011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(24),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(24),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010000011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010000011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(26),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010000011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010000011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(28),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(28),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010000011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010100111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010000011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010000011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101001010000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101001010000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(43),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010011010010101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010100111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101001010000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010000011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010000011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(21),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(21),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010000011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(22),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(22),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010000011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(35),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101001010000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101001010000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101001010000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(38));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101001010000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101001010000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101001010000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(40),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(40));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101001010000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101001010000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(46),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010000011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010011010010101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101001010000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(54));
GRLFPC2_0_COMB_UN1_R_A_RS1_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001011110010")
port map (
combout => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\,
dataa => \GRLFPC2_0.R.A.RS1\(0),
datab => \GRLFPC2_0.R.A.RS1D\,
datac => \GRLFPC2_0.COMB.UN1_FPCI_3_1_X\,
datad => \GRLFPC2_0.COMB.UN4_LOCK_0\);
GRLFPC2_0_COMB_RS2D_1_IV_0_O2_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100001101100000")
port map (
combout => \GRLFPC2_0.COMB.RS2D_1_IV_0_O2_0\,
dataa => N_69,
datab => N_76,
datac => N_66,
datad => N_64);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(46),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(43),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(45),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(50));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(35));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(35));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110110001101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_T_3_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011001110110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_T_3\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(377),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.SELECTQUOBITS.NOTDIVC\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.SELECTQUOBITS.NOTDIVC\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD57\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(20),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(21),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(20),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(28),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_3_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111100001110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3_A\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_3_A_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3_A\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(256),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_235_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111000010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_235__G0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(235),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0\(235),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M2_0\);
GRLFPC2_0_COMB_UN1_FPCI_4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001011110010")
port map (
combout => \GRLFPC2_0.COMB.UN1_FPCI_4\,
dataa => \GRLFPC2_0.R.A.RS2\(0),
datab => \GRLFPC2_0.R.A.RS2D\,
datac => \GRLFPC2_0.COMB.UN1_FPCI_3_1_X\,
datad => \GRLFPC2_0.COMB.UN4_LOCK_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100111011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPAREGLOADEN_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datab => \GRLFPC2_0.FPI.LDOP_REP0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.WQSCTRL\(68),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN53_SCTRL_NEW: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.UN53_SCTRL_NEW\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.U_RDN_1\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010100111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(8),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010000011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101001010000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101001010000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101001010000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(50));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_6\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101001010000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101001010000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(45),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(45));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_UN3_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.UN3_TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.TEMP_25_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.TEMP2_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.UN4_TEMP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN10_S_MOV\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_236_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111000010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_236__G0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(236),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0\(236),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M2_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_NORMDETECT_NOTSLFROMNORM_19_3_0__M2\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010001110100011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19_3_0_.M2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M14\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_NORMDETECT_NOTSLFROMNORM_19_3_0__M3\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010001110100011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19_3_0_.M3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M14\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_NORMDETECT_NOTSLFROMNORM_19_3_0__M4\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010001110100011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.NORMDETECT.NOTSLFROMNORM_19_3_0_.M4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M14\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110101001101010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.EXPYBUS_0\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110101001101010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.EXPYBUS_0\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110101001101010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.EXPYBUS_0\(7));
GRLFPC2_0_COMB_UN3_IUEXEC_RNI88491: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101111")
port map (
combout => \GRLFPC2_0.COMB.FPOP_0_0_O2\,
dataa => N_89,
datab => N_90,
datac => \GRLFPC2_0.COMB.FPOP_0_0_O2_0_2\,
datad => \GRLFPC2_0.COMB.UN3_IUEXEC\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN30_CONDITIONAL_M5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111100010101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN30_CONDITIONAL_M5\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN30_CONDITIONAL_M2_E_4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN30_CONDITIONAL_M2_E_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN30_CONDITIONAL_M5_A\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN30_CONDITIONAL_M5_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010101010111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN30_CONDITIONAL_M5_A\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD9\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD10\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_14_RNIS66H_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110010100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_9__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_10_1\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_9_0_A2\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_14\(34));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CONDMUXMULXFF.UN4_NOTSQRTLFTCC\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_1_RNI8DSK_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A3\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_14_2\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_14_1\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_1\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_0_RNIB57H_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_17__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_16_1\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_O28_5\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_2_0_A2\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_2\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_O2\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_14_0_A2\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010011110100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_1_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_6_I_O2\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7_2\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_11_0_A2\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_0_I_O2\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101011000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_4859_A2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_36\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_18_2\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_26_2\(60));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_13_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8466_I_I_I_X2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_2\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_8\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_9_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_1\,
dataa => N_32980_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_22_1\(58),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_15\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101011000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_6_0\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_4859_A2_1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_1_0_A2\(62),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_26_2\(60));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2_0\,
dataa => N_34381_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_4785_A2_2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\(58),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(50));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A13_1\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_13_1\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_2\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_11_0\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_1\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_18\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_2\(25),
datab => N_28709_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_12_0\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_9\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN1_S_DYADIC_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_2\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_2\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_39__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_9_0_A2\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_14_1\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(38));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110010100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_16_0\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_15_0\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_16_1\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_10_1\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_5\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_14_2\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_10\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2_2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_7_2\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_2\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_10\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_0\,
dataa => N_33495_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_4_0\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_14\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_0_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_0\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_1_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8577_I_0_A2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_12\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_6_1\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_10_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_6\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_0_2\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_2\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_12\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_13_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A13_0\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_2\(57),
datac => N_28871_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_4\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_18_3\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_17\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_16_1\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_2_1\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_19\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_7_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_2_4\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_4\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_5_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_3_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_0_2\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_11\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_6_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_13_1\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_1\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_9\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_6\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_6_1\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_1\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A15_1\(18),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_14_2\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_10\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_1_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_16_1\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_6_1\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_22\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_4\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_3\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_0_7_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_7\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A28_1\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_O28_1\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_2\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_2\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_0_6_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011110111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_6\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_11_0\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\(58),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_9\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_0_1_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_1\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_9_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_2\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_3\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_0_0_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011101110111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_0\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_6_0\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_O28_5\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_14_1\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_9_1\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_9_0\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_5\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_11_0\(18),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_11_2\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_13_1\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_5\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_16_2\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_14_3\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_12\(60));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_4_RNIUTQG_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_3\,
dataa => N_33495_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_4\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_4_RNI03PQ1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0_1\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_4\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_6_RNINRLB_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_0\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_9_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_14_1\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_6\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101110000001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_8\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O18_4\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_7_0\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_10_1\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_5\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_5\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_8\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_6\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_13_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_13_2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A26_1\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_5\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_2\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_2_0\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_5_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_14\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_17_1_0\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0_1\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_6\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_10_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_16_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_O28_5\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_5_1\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_10\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_11_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_M2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_O28_5\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_5\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_9_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_4_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_3\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_2\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_1_9_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011101110111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_9\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_10_1\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_17_2\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_1_8_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001101011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_8\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_X2_2\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_2\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_16_2\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_1\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_1_6_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_6\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_20_2\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_2_1\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A26_1\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_3\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_1_5_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011101110111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_5\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_9_0\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_9_1\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_4\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A21_1\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_3_0_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_3_0\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_11_0\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_5_0\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_1_2_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_2\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80),
datab => N_33495_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_15_3\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_6\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_1_1_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111100000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_1\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_2\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_2_1\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_13\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_1_0_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_0\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_1_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_11_2\(5),
datac => N_29496_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_0\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_13_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_10\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_2\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_2_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_14_1\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_11\(60));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_10_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_8\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_2\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_O30_7\(60),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_8\(60));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101000110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_5\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_2_0\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_2\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_10_0\(60),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_27_1\(60));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_1_1\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O2\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_16_1\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_4\(60));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_5_0\(60),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_17\(60));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_1_1_0\(62),
datab => N_33227_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_I_X2\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_7\(62));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_5_1\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_7\(62));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A29_RNID639_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_8_1\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1_A2_1_1\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A30_22_RNIDNQB_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_6\,
dataa => N_33157_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_8_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_22\(60));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_2_2_RNI5QCE_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_19__G2_4\,
dataa => N_32980_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_3_1\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_2_2\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_21\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_11\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O25\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_9\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_0\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O2\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_20\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_16_1\(51),
datab => N_28709_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O2\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_0\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_13_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_2_1\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O2\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_4\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_6\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_8_1\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_15\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_9_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A3\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_1_1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_2_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_10\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_1_1\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_20_0\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_12\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_4_1\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O18_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_10_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101011000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_5\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_17_1\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_10_0\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_11\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_17_0\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_11_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_14_0\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O21\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_21\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_9_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_22_1\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O21\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_4\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_1_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_13\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_15__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_14_2\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_27\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A15_0\(18),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_14_0\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_17_1\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_26_2\(60));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_9\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_1\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_2\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_6_1\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_19\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_8\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A13_1\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_21_1\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_2\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_10_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_8_1\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_16_1\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_12_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_13\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_16_1\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_20_1_0\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_12\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A13_1\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_14\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_2_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_9_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_8\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_8_A\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_12_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011011111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_8_A\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X3\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_10_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_5\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_1\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_21\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_13_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_10_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_9\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_1\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0_1\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_4\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A15_1\(18),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_10_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_5_1\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_7\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000111110001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_0\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_2_3\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_0_I_O2\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_26_2\(60));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_7_2\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_4\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_13_1\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_1\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_1\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_9_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101011000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_10_0\(34),
datab => N_33157_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_9_0\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A22_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_6_2\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_13_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_12_0\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O2\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_5\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110010100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_1_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_2_1\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_8_0\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_0_2\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_12_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_3_1\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_15_1\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_23\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_I_A26_1\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_38\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_7_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_5_3\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_37\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_11_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_12_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_30\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010100001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_1_A\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_10_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001011000000110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2_1_A\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83),
datad => N_32980_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_6_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_0\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(58),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_4\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_2\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_0\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_12_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_7\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_1_1\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_21_2\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_13\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2_1\,
dataa => N_33157_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_4\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_5_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_24\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_1_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_O2\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2\(42));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_ENTRYPOINT_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.ENTRYPOINT_1\,
dataa => N_33495_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_1_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8577_I_0_A2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN10_S_MOV\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_ENTRYPOINT_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.ENTRYPOINT_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_7_1\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN1_S_DYADIC_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.S_CMP\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_12_2_RNILURA_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110010100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A19_1\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_12_2\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_7_2\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_2_0_A2\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_10_1_0_A2_RNIN57G_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000111110001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_10_1_0_A2\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0_1\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_6_I_O2\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_17_2\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_2_0_O2_0_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_2_0_O2_0\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_0\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_O2\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_2_A2_1\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_0_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_0\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_16_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_8_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_11_0_A2\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_0_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100011111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_44__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0_0\(43),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_4_2\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_1_0_A2\(62),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_O2\(25));
GRLFPC2_0_R_A_LD_RNO_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000000000000")
port map (
combout => \GRLFPC2_0.R.A.LD_0_0_G1_3\,
dataa => N_76,
datab => N_77,
datac => N_88,
datad => \GRLFPC2_0.R.A.LD_0_0_G1_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0_0_A2_RNIV8VF_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_12__G2_2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_4_1\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_26_2\(60),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_0_0_A2\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_0_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_0\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(42));
GRLFPC2_0_COMB_UN6_IUEXEC_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100010")
port map (
combout => \GRLFPC2_0.COMB.UN6_IUEXEC_1\,
dataa => \GRLFPC2_0.R.MK.BUSY2_RET_1\,
datab => \GRLFPC2_0.R.MK.BUSY2_RET\,
datac => \GRLFPC2_0.R.MK.BUSY_RET_4\,
datad => \GRLFPC2_0.COMB.UN6_IUEXEC_1_A\);
GRLFPC2_0_COMB_UN6_IUEXEC_1_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.COMB.UN6_IUEXEC_1_A\,
dataa => \GRLFPC2_0.R.MK.BUSY_RET_5\,
datab => \GRLFPC2_0.R.MK.BUSY_RET_2\,
datac => \GRLFPC2_0.R.MK.BUSY_RET_3\,
datad => \GRLFPC2_0.R.MK.BUSY_RET\);
GRLFPC2_0_N_939_I_I_A2_1_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001110000000000")
port map (
combout => \GRLFPC2_0.N_939_I_I_A2_1_0\,
dataa => N_77,
datab => N_87,
datac => N_80,
datad => N_78);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN3_NOTAZERODENORM_RNI989G: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010100010101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_0\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN3_NOTAZERODENORM\);
GRLFPC2_0_R_I_RDD_RNO_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.R.I.RDD_0_0_G1_0_8238_I_A3_1\,
dataa => \GRLFPC2_0.R.A.MOV_RET\(15),
datab => \GRLFPC2_0.R.A.MOV_RET\(12),
datac => \GRLFPC2_0.RS2_0_SQMUXA_3\,
datad => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_11\);
GRLFPC2_0_COMB_ANNULFPU_1_U_0_O2_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101011000000")
port map (
combout => \GRLFPC2_0.COMB.ANNULFPU_1_U_0_O2_0\,
dataa => \GRLFPC2_0.COMB.UN1_FPCI_2_X\,
datab => \GRLFPC2_0.COMB.UN1_FPCI_X\,
datac => \GRLFPC2_0.R.X.FPOP\,
datad => \GRLFPC2_0.R.E.FPOP\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_5\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_13_1\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_5_TZ\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_5_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_0_S\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_OPREXC_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_4\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_5\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN3_NOTBZERODENORM\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTDECODEDUNIMP_A_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010100000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN1_S\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN6_S\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_13_2\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_8_0\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O25\(27));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN2_INEXACT: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN2_INEXACT\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN2_INEXACT_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.NOTAM2\);
GRLFPC2_0_COMB_UN8_CCV: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000111")
port map (
combout => CPO_CCVZ,
dataa => N_352,
datab => \GRLFPC2_0.R.X.FPOP\,
datac => \GRLFPC2_0.COMB.UN8_CCV_0\,
datad => \GRLFPC2_0.COMB.UN8_CCV_1\);
GRLFPC2_0_COMB_UN1_MEXC_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111000000000000")
port map (
combout => \GRLFPC2_0.COMB.UN1_MEXC_1\,
dataa => \GRLFPC2_0.R.FSR.TEM\(4),
datab => \GRLFPC2_0.R.I.EXC\(4),
datac => \GRLFPC2_0.COMB.UN1_MEXC_1_0\,
datad => \GRLFPC2_0.COMB.UN1_MEXC_1_1\);
GRLFPC2_0_COMB_V_A_AFSR_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.COMB.V.A.AFSR_1\,
dataa => \GRLFPC2_0.COMB.V.A.AFSR_1_1_0\,
datab => \GRLFPC2_0.N_782\,
datac => \GRLFPC2_0.COMB.V.A.AFSR_1_2\,
datad => \GRLFPC2_0.COMB.UN4_LOCK_0\);
GRLFPC2_0_COMB_V_A_AFQ_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101000000000000")
port map (
combout => \GRLFPC2_0.COMB.V.A.AFQ_1\,
dataa => \GRLFPC2_0.R.A.SEQERR_RET_4\(0),
datab => \GRLFPC2_0.R.A.SEQERR_RET_4\(1),
datac => \GRLFPC2_0.COMB.V.A.AFQ_1_6\,
datad => \GRLFPC2_0.COMB.V.A.AFQ_1_10\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_0\,
datac => \GRLFPC2_0.FPI.LDOP_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP0\);
GRLFPC2_0_COMB_UN2_HOLDN_0_A2_13: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_13\,
dataa => \GRLFPC2_0.COMB.UN3_HOLDN_X\,
datab => \GRLFPC2_0.R.A.FPOP\,
datac => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_13_3\,
datad => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_13_4\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CHECKOVANDDENORM_UN13_NOTPOSSIBLEOV: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD51\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD52\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_4\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN26_NOTBINFNAN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN26_NOTBINFNAN\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN8_NOTBINFNAN\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN26_NOTBINFNAN_4\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN26_NOTBINFNAN_5\);
GRLFPC2_0_COMB_FPDECODE_RS1D5_0_A2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.COMB.FPDECODE.RS1D5_0_A2\,
dataa => N_66,
datab => N_65,
datac => \GRLFPC2_0.COMB.FPDECODE.RS1D5_0_A2_0\,
datad => \GRLFPC2_0.RS1V_0_SQMUXA_1_0_A2_2_X\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_26_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_26\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_16_2\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_14_1\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79),
datab => N_33157_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_8_2\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_5_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_5\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_0_A2\(46),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_3_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_3\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_1\(5),
datab => N_33227_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_13_2\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_14_1\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A7_3_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_3\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_13_0\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A7_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A7\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O7_2\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_4_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_4\(32),
dataa => N_28709_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_2\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_4_1\(50),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_7_1\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_2_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_2\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_1_1\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O20_3\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_1_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_1\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_13_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_1_1\(62),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_2_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A6_3_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A6_3\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O6\(30),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_14_1\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A6_2_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A6_2\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_9_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_13_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A6_2_1\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_17_1_I_O2\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_5_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_2_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_2\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_12_0_A2\(62));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_1_A2_0_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1_A2_0\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8466_I_I_I_X2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_7_1\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_25_1\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_1_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_1\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_3\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_25_1\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0_0\(12),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A16_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A16\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_1\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_5_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_12_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_0_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_0\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_1_1\(62),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_1\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A23_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7_1\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_1_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_1\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_7\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_0_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_0\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_0_2\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_13_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_2\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_7_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_7\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_10_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O29_1_0\(58),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_2_2\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_10_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_10\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8466_I_I_I_X2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_0_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_0\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_4_1\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_8_1\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_12_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_3_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_3\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_5\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0_1\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_0_A28_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_A28\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A7_1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A2_7\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A28_0_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_0\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_0_S\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_3_1\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_1\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A26_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A26\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O26_9\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A26_1\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_0_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_0\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_2\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O26_8\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_1_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_1\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11_1\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_5_1\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_3_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_3\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_7_1\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O26_5\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_20_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_20\(53),
dataa => NN_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_0\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O2\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_21_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_21\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_9\(53),
datac => N_33495_1,
datad => N_29496_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_29_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_29\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_0\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_2_1\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_0_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_0\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_1_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_0_0\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_4\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_1_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_1\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_16_2\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_1\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_1_2\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_O27_4\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_6_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_6\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_6_0\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_7_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_2\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A25_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A25\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_7\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A19_1\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A25_1\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_1_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_1\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_1\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_1\(59),
datad => N_34483_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_2_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_2\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A19_1\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_1_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_2_0\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A24_7_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_7\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_1_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_7_0\(11),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_0_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_0\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_18_1_0\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O2\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A27_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A27\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_1\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(13),
datad => N_34483_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_0_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_0\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_1\(59),
datab => N_33157_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_5\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A19_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A19\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A19_2\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_4\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A13_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A13\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A13_0\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_1\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8577_I_0_A2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A21_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A21\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN1_S_DYADIC_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A21_1\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_0_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_4_2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0_0\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0_1\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_5_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_5\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_M21\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_1_1\(62),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_6_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_6\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_1\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_13_1\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_1\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A28_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A28\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A28_1\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_M2_0\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_1_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_1\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_1_1\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O28_5\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O2\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_I_A26_3_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_3\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A13_1\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_O2_2\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O25\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_1_0\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_12_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_0_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_0\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_0_2\(36),
datac => N_28709_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0_1\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_2_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_2\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_2_0\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_5\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_12_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_3_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_3\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_3_1\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_9_0\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_2\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A21_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A21\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A21_2\(51),
datab => N_33495_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_5_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_13_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_6_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_6\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_18\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_12_1\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A7_0_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_0\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_0_1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A7_1_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_1\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_5\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A3\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_19\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_0_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_2\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_14_2\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_12_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_1_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_1\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O18_6\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O13_0\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_2_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_2\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_3_1\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_2_1\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A25_1\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_5_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_5\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(59),
datab => N_32980_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_5_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_2\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_2\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_2_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_8_1\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_1_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_1\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_4_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_1_1\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_1_2\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_13_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_7_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_7\(48),
dataa => N_28709_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_7_2\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_5_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_4_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A3\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN1_S_DYADIC_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_1\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A30_1_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_1\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_1_0\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_5_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_1_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_1\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_1_0\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_6\(13),
datad => N_34483_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_3_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_3\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_1_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_3_1\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_6_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_6\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_7_1\(34),
datac => N_33157_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_8_1\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_5_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_5\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_5_0\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_0_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_0\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_7_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_O27_2\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_6_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_6\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_7_1\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_6_0\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_3_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_3\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_10_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_3_1\(58),
datad => N_28871_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_5_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_5\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_5_0\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_13_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_3_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_3\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_2\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_1_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_1\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_3_1\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_1_1\(19),
datad => N_34072_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_3_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_1_1\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_1\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_12_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_2_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_2\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_1_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_10_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_19\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_2_0\(35),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A7_0_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_0\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_5_1\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_0_1\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_4_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_4\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_10_1\(11));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP2_0_RNI61T11: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.TEMP_25\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.TEMP_25_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.TEMP2_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN10_S_MOV\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A18_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A18\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_16_1\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_5\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O18_0\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010011000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_8645\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A3\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_8645_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_7_0\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_9_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010111000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_0_2\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(58),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_10_1\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_12_2\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2_3_TZ\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_9_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O18_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_3_1_0\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_12_RNIGK6G_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_14_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_12\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_0_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110000001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_0\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_0_0\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O2\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_2\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_YY_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101000110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_YY\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_YY_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101000110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_YY\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_YY_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101000110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_YY\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_YY_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101000110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_YY\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_9_TZ_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001100110011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_9_TZ\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_22_0\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_14_2\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111000011110100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2_5_TZ\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_1_0_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O13_0\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_8_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => N_34381_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11_2\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_16_1\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_2_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_17_1_I_O2\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_16_1\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_O2\(25));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SIGNRESULT: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110000001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.SIGNRESULT\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(23),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SFTLFT.UN1_GRFPUS\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN20_ZERO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111001111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN23_EXPXBUS_10_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001100110011001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.UN23_EXPXBUS_10_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(10));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN5_SHDVAR: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111011101110111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN5_SHDVAR\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_0\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_0\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.EXPYBUS\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.EXPYBUS\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_RNIO9A6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_RNIF0H2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_3_RNI4R37: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_2_RNI8RN3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_1_RNIPP32: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_RNIKB7E: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_RNIB2EA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_2_RNI5VSA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_2_RNIAVG7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_1_RNIEV44: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_3_RNI61V1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_2_RNIKVO8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_RNINLS6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_3_RNIQPS3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_2_RNIBO82: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_RNILMD9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN50_ZERO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111001111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_3_RNI9KV7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_1_RNICKJ4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_2_RNIIK79: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_1_RNI7LN3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_2_RNIDLB8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_2_RNI3KB3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_1_RNIODUC: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_3_RNIEGQ4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_3_RNIDGQ4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_1_RNI7QV7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_1_RNI8P06: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_1_RNIDPK2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_3_RNIKP87: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_3_RNIPPS3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_2_RNIAO82: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_2_RNIFOS6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_RNIBDK5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_2_RNIPO48: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_RNIPQ16: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_RNI7864: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_3_RNI5KB3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_3_RNIAKV7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_1_RNIDKJ4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_1_RNIIK79: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_1_RNINKR5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_RNIADB3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_RNIKC14: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_2_RNI61V1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_1_RNIAGQ4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_3_RNIBGQ4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_3_RNIAGQ4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_2_RNI3QB3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_3_RNIOKR5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_2_RNISKFA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_RNI04I7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_1_RNI5LN3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_3_RNIDLB8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_1_RNIGLV4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_1_RNI7GQ4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_1_RNI6GQ4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_1_RNIOE52: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_3_RNIVEP6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_1_RNI2FD3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_3_RNI9F18: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_1_RNICFL4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_RNI14I7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_3_RNILE2C: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_2_RNIEV44: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_2_RNIJVO8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_RNIDIJ4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_RNIT5N6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_1_RNIEUC8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_3_RNILU05: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_2_RNI8VG7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_RNIU464: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_RNILRC8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_3_RNIOVC5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_RNIS5N6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_2_RNIEUC8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_2_RNISFH2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_1_RNI0G57: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_1_RNI56S: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_3_RNIC6G5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_RNI5PA1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_RNI3ABB: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_1_RNIUU86: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_1_RNI3VSA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_RNI8EV7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_2_RNI9L05: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_3_RNISJC3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_2_RNICLB8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_3_RNIILV4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_RNI2ABB: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_3_RNIVU86: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_3_RNI4VSA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_RNIAJ47: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_RNI1ABB: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_RNIO0I7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_1_RNIKKGA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_3_RNIRK47: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_RNIGQP3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_1_RNI3LC8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_2_RNIIQ79: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_RNIQQ16: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_3_RNI5PC9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_1_RNIOEM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_1_RNIAD27: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_1_RNIFDMB: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_2_RNILDA8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_2_RNIQDUC: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_3_RNI0EI9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_2_RNI4E6E: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_1_RNI8EQA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_2_RNIEEE7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_RNIMAMB: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_1_RNINEM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_RNITK0A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_1_RNIUPN6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_2_RNIDQJ4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_3_RNIOQR5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_3_RNIGEE7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_3_RNIMOG3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_3_RNIRO48: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_1_RNIMFT5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_2_RNI6GP3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_2_RNIOE52: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_RNI2DA9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_3_RNI3FD3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_3_RNI8F18: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_2_RNICFL4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_3_RNIIF99: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_2_RNIMFT5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_3_RNI8LN3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_1_RNI15G: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_1_RNI6545: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_3_RNID5O1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_RNIQG28: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_3_RNIS5K7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_2_RNI0684: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_RNID245: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_RNI4PA1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_1_RNIC1V1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_RNIPFRA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_RNIG627: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_1_RNI7EQA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_2_RNIDEE7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_1_RNIIE2C: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_2_RNIOEM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_RNI3LJA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_1_RNIK9H8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_2_RNI0K08: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_2_RNI5KK4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_3_RNIBK89: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_UN120_TEMP_0_RNIFMDJ: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.UN123_TEMP_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.UN120_TEMP_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_UN123_TEMP_0_RNI3V0K: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.UN126_TEMP_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.UN123_TEMP_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_UN126_TEMP_0_RNIN7KK: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.UN129_TEMP_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.UN126_TEMP_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_UN132_TEMP_0_RNIIICL: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.UN129_TEMP_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.UN132_TEMP_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_RNIMBT: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_RNIOC14: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_1_RNI91V1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_2_RNIM503: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_RNIPC14: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_2_RNIEGQ4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_3_RNI6GR4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_2_RNI4GR4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_2_RNI3LC8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_3_RNI9L05: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_2_RNI6GR4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_1_RNIG9H8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_2_RNIG9H8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_2_RNI3GR4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_2_RNI2GR4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_2_RNI1GR4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_1_RNIVFR4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_RNIMC14: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_RNILC14: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_CIN_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.CIN_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_1_RNI2PC9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_RNI78F6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_RNIV752: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_RNI5NN6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_2_RNIUFH2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_1_RNI2G57: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_1_RNIOVC5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_3_RNICUO3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_2_RNIGUC8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_RNIDM35: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_3_RNI0FP6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_1_RNIJ9H8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_3_RNIUFH2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_1_RNI1G57: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_RNI0LJA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_3_RNIJ9H8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_RNISKJA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO_REP2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_1_RNI3QB3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_1_RNI8QV7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_2_RNIEQJ4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_RNI0J32: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_2_RNIOQR5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_RNIE0H2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_2_RNI7RN3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_3_RNIQP32: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_RNI3O89: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_V\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_RNICJ47: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_V\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_2_RNI4FD3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_2_RNI9F18: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_3_RNIFFL4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_3_RNIGGQ4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_V\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN50_ZERO_REP2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_RNIT203: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_2_RNIJF99: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_3_RNIPFT5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_1_RNI6GP3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_V\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC2_0_COMB_RDD_1_M14_0_O2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111100100000")
port map (
combout => \GRLFPC2_0.COMB.RDD_1.M14_0_O2\,
dataa => N_65,
datab => N_64,
datac => N_67,
datad => N_68);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_114_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(114),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(114),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(114),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_2_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100000001111")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_2\(3),
dataa => \GRLFPC2_0.R.I.EXC\(3),
datab => \GRLFPC2_0.R.FSR.TEM\(3),
datac => \GRLFPC2_0.COMB.V.FSR.CEXC_1_2_A_X\(3),
datad => \GRLFPC2_0.COMB.V.FSR.CEXC_1_SN_M2\);
GRLFPC2_0_COMB_RDD_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110011001100")
port map (
combout => \GRLFPC2_0.COMB.RDD_2\,
dataa => \GRLFPC2_0.R.X.RDD\,
datab => \GRLFPC2_0.R.I.RDD\,
datac => \GRLFPC2_0.R.I.RDD_0_0_G1_0_8238_I_O4\,
datad => \GRLFPC2_0.COMB.UN1_R.I.V_0\);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_2_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100000001111")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_2\(1),
dataa => \GRLFPC2_0.R.I.EXC\(1),
datab => \GRLFPC2_0.R.FSR.TEM\(1),
datac => \GRLFPC2_0.COMB.V.FSR.CEXC_1_2_A_X\(1),
datad => \GRLFPC2_0.COMB.V.FSR.CEXC_1_SN_M2\);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_2_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100000001111")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_2\(4),
dataa => \GRLFPC2_0.R.I.EXC\(4),
datab => \GRLFPC2_0.R.FSR.TEM\(4),
datac => \GRLFPC2_0.COMB.V.FSR.CEXC_1_2_A_X\(4),
datad => \GRLFPC2_0.COMB.V.FSR.CEXC_1_SN_M2\);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_2_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100000001111")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_2\(2),
dataa => \GRLFPC2_0.R.I.EXC\(2),
datab => \GRLFPC2_0.R.FSR.TEM\(2),
datac => \GRLFPC2_0.COMB.V.FSR.CEXC_1_2_A_X\(2),
datad => \GRLFPC2_0.COMB.V.FSR.CEXC_1_SN_M2\);
\GRLFPC2_0_COMB_V_FSR_CEXC_1_2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100000001111")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_2\(0),
dataa => \GRLFPC2_0.R.I.EXC\(0),
datab => \GRLFPC2_0.R.FSR.TEM\(0),
datac => \GRLFPC2_0.COMB.V.FSR.CEXC_1_2_A_X\(0),
datad => \GRLFPC2_0.COMB.V.FSR.CEXC_1_SN_M2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(45),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(180),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(46),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(20));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100011111011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011001011111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(24),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0_A\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_A_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010110011101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0_A\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0_A\(25));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_A_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010110011101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0_A\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(26),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(21),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(22),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(28),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(26),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0_A\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_A_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001100101011101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0_A\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(29),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(14));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010011111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(22),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(24),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0_A\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_A_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010110011101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0_A\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(23),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(25));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010011111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0_A\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_A_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010110011101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0_A\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(24),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(50));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(40),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(40));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(46),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(201),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(38));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(35),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0_A\(35));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_A_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010110011101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0_A\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(38));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000111101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000111101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111001001110010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3_A\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_A_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3_A\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111001001110010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3_A\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_A_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3_A\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_3_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.U_RDN_1\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(35));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(45),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(43),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0_A\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_A_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001100101011101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0_A\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(30),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(25));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(40),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(40));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111011100001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3_A\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_A_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001101100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3_A\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(21),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(22),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(20));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(22),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(28),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(50));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_3_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_2\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_1\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_3_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2_1\(9),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3_A\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_3_A_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3_A\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(241),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(254),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_0\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_0\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_173_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_173__G0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(173),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14_142_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011110010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_14\(142),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(144),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLCREGXZ.UN11_INFORCREGSN\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_RNIGPS6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRTOSTICKY\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TEMP\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD10\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD11\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN12_SRTOSTICKY_3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(183),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(48));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN35_ZERO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111001111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN5_ZERO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_A\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_UN5_ZERO_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_A\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(20));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(14));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3_A\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_A_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3_A\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(50),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3_A\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_A_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3_A\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_3_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_3\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN1_TEMP\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW\(77),
datad => \GRLFPC2_0.FPI.LDOP_REP1\);
GRLFPC2_0_V_FSR_FTT_1_SQMUXA_3_0_RNIRQVN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101011111010")
port map (
combout => \GRLFPC2_0.UN1_FPCI_21\,
dataa => \GRLFPC2_0.COMB.UN1_FPCI_X\,
datab => \GRLFPC2_0.R.X.AFQ\,
datac => \GRLFPC2_0.V.FSR.FTT_1_SQMUXA_3_0\,
datad => \GRLFPC2_0.N_1213_I_0_O2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(38));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M14_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M14\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M14S2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M14_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M14\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M14S2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M14_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M14\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13_0\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M11S4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M14S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_3_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_2\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_1\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_3_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_2\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_1\(7));
GRLFPC2_0_COMB_FPDECODE_FPOP3_0_A2_1_X_RNI80AG: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.COMB.RS1_1_SN_M2_I_A2\,
dataa => N_88,
datab => N_87,
datac => \GRLFPC2_0.COMB.FPDECODE.ST_0_A2_0_A2_0_X\,
datad => \GRLFPC2_0.COMB.FPDECODE.FPOP3_0_A2_1_X\);
GRLFPC2_0_COMB_FPDECODE_FPOP3_0_A2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.COMB.FPDECODE.FPOP3_0_A2\,
dataa => N_80,
datab => N_77,
datac => N_76,
datad => \GRLFPC2_0.COMB.FPDECODE.ST_0_A2_0_A2_0_X\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_7_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010110011101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_7_A\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SFTLFT.AREGXORBREG_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD12\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSRRES_0_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSRRES_0\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(20));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_2_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_2\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_34_2\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_6_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_6\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_36\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_14_1\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_4_0_A2_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_4_0_A2\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_16_2\(6),
datac => N_34381_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000011100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN1_S_DYADIC_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_35\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_10_1\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000110100001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_35\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_O2\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_1_A2_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1_A2\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_2\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_2_0_A2\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1_A2_3\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0_A2_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_0_A2\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_16_2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O18_4\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_O28_5\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0_A2_0_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_0_A2_0\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_16_2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A26_1\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_7_2\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_12\(60));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100011111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_2_0_A2\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_26_2\(60),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_17\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0_0_O2_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101011000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_0_0_O2\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_8_1\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN1_S_DYADIC_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_13_2\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_2_1\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O6_3_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111000011110010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O6_3\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_9_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_2_1\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_10_2\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_14_1\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O29_6_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110010100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O29_6\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_10_1\(4),
datab => N_33157_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_1_2\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O23_6_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011000111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_6\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_M2_0_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010100011111101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_M2_0\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_O2_1_0\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_13_1\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_O2_3\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O7_1_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000111110001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O7_1\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A19_1\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A3_3_2\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_0\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_2_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_2\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_8_1\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O13_0\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_3_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_3\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_8_1\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O13_0\(0));
GRLFPC2_0_R_A_LD_RNO_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC2_0.R.A.LD_0_0_G1_0\,
dataa => N_81,
datab => N_79,
datac => N_92,
datad => \GRLFPC2_0.N_939_I_I_2_0_X\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A7_0_1_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_0_1\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_4_1\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_0_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101000001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0_0\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_2_2_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_2_2\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_5_1\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_9_3_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_9_3\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_8_1\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_9_1\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A7_0_1_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_0_1\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_2\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_1_1_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_1_1\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_0_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0_0\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8466_I_I_I_X2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_0_1_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_0_1\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_5_0_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010011100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_5_0\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_5_1\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_10_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_10_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_10_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_16_1_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001011100010111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_16_1\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_5_2_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_5_2\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_1\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A14_2_3_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_2_3\(62),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => N_33227_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_1\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A6_2_1_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A6_2_1\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_3_1_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_3_1\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_0\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_1_0_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_1_0\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8466_I_I_I_X2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_0_1_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_0_1\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_0\(34));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN11_INEXACT_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN11_INEXACT_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(39),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(40),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_6_1_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_6_1\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_7_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_2_1_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_2_1\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_0_1_0_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0_1_0\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A15_1\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_16_1_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_16_1\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79),
datad => N_33495_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_2_1_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_2_1\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A3\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRLEN_RNO_8_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_13__G2_3_TZ_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_2_1\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_1\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_7_1_0_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_7_1_0\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83),
datad => N_32980_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_4_1_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_4_1\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_2\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_4_1_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_4_1\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_1\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_8_1_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_8_1\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_9_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_9_1_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_9_1\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_11_2\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_24_1_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_24_1\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_2_1\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_10_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A24_8_1_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_8_1\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_3\(51));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_24: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_24\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_20\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_23: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_23\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_9\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_19\);
GRLFPC2_0_COMB_ANNULFPU_1_U_0_O2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110010100000")
port map (
combout => \GRLFPC2_0.COMB.ANNULFPU_1_U_0_O2_1\,
dataa => \GRLFPC2_0.COMB.UN1_FPCI_1_X\,
datab => \GRLFPC2_0.COMB.UN3_HOLDN_X\,
datac => \GRLFPC2_0.R.M.FPOP\,
datad => \GRLFPC2_0.R.A.FPOP\);
GRLFPC2_0_COMB_V_A_AFQ_1_10: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.COMB.V.A.AFQ_1_10\,
dataa => \GRLFPC2_0.R.A.AFQ_RET_5\,
datab => \GRLFPC2_0.R.A.ST_RET_2\(0),
datac => \GRLFPC2_0.COMB.V.A.AFQ_1_4\,
datad => \GRLFPC2_0.COMB.V.A.AFQ_1_7\);
GRLFPC2_0_R_E_SEQERR_RNO_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.COMB.SEQERR.UN3_QNE_3\,
dataa => \GRLFPC2_0.R.A.MOV_RET\(12),
datab => \GRLFPC2_0.R.A.MOV_RET\(13),
datac => \GRLFPC2_0.COMB.QNE2_0\,
datad => \GRLFPC2_0.COMB.V.A.AFSR_1_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN2_INEXACT_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN2_INEXACT_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(39),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(40),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(10));
GRLFPC2_0_RIN_MK_LDOP_9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC2_0.RIN.MK.LDOP_9\,
dataa => \GRLFPC2_0.R.MK.LDOP_RET_1\(3),
datab => \GRLFPC2_0.R.MK.LDOP_RET_1\(0),
datac => \GRLFPC2_0.RIN.MK.LDOP_6\);
GRLFPC2_0_RS1V_0_SQMUXA_1_0_A2_0_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.RS1V_0_SQMUXA_1_0_A2_0_1\,
dataa => N_65,
datab => N_64,
datac => \GRLFPC2_0.RS1V_0_SQMUXA_1_0_A2_3_X\,
datad => \GRLFPC2_0.RS1V_0_SQMUXA_1_0_A2_1_X\);
GRLFPC2_0_COMB_RDD_1_M14_0_A2_1_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC2_0.COMB.RDD_1.M14_0_A2_1_1\,
dataa => N_87,
datab => N_80,
datac => N_88,
datad => N_78);
GRLFPC2_0_RS1D_CNST_0_A3_0_A2_0_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC2_0.RS1D_CNST_0_A3_0_A2_0_0\,
dataa => N_80,
datab => N_77,
datac => N_87,
datad => \GRLFPC2_0.COMB.FPDECODE.RS1D5_0_A2_0\);
GRLFPC2_0_RS1V_0_SQMUXA_1_0_A2_2_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110000000000000")
port map (
combout => \GRLFPC2_0.RS1V_0_SQMUXA_1_0_A2_2_0\,
dataa => N_62,
datab => N_63,
datac => \GRLFPC2_0.RS1V_0_SQMUXA_1_0_A2_1_X\,
datad => \GRLFPC2_0.RS1V_0_SQMUXA_1_0_A2_2_X\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_3_1_0_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_3_1_0\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O18_4\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_11_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010101000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_6\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_3_1\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_1\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O25\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(33));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN17_SHDVAR: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR_A\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN17_SHDVAR_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101010100000011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR_A\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_U_RDN_1_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.U_RDN_1\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.UN6_U_RDN\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_S_CMP: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.S_CMP\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_1_1\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_10_1\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(52));
GRLFPC2_0_COMB_UN2_HOLDN_0_A2_11: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011100000000")
port map (
combout => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_11\,
dataa => \GRLFPC2_0.R.A.MOV_RET\(4),
datab => \GRLFPC2_0.R.A.MOV_RET\(5),
datac => \GRLFPC2_0.R.A.MOV_RET\(11),
datad => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_11_0\);
GRLFPC2_0_COMB_UN4_LOCK_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011110010")
port map (
combout => \GRLFPC2_0.COMB.UN4_LOCK_0\,
dataa => \GRLFPC2_0.R.A.SEQERR_RET_4\(0),
datab => \GRLFPC2_0.R.A.SEQERR_RET_4\(1),
datac => \GRLFPC2_0.COMB.UN4_LOCK_0_2\);
\GRLFPC2_0_R_I_EXC_RNO_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC2_0.R.I.EXC_2_0_3__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(38),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(40),
datad => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2\);
\GRLFPC2_0_R_I_EXC_RNO_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000010000")
port map (
combout => \GRLFPC2_0.R.I.EXC_2_0_1__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(40),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DECODESTATUS.UN7_STATUS\,
datad => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2\);
GRLFPC2_0_R_MK_BUSY_RET_4_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.R.MK.BUSY_RET_4_0_0_A2_0_G0\,
dataa => \GRLFPC2_0.R.MK.RST_RET_3\,
datab => \GRLFPC2_0.R.MK.RST_RET_2\,
datac => \GRLFPC2_0.R.MK.BUSY_RET_4_0_0_A2_0_G0_2\,
datad => \GRLFPC2_0.R.MK.BUSY_RET_3_0_0_A2_X\);
GRLFPC2_0_COMB_V_MK_RST_1_0_A2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.COMB.V.MK.RST_1_0_A2\,
dataa => \GRLFPC2_0.R.MK.HOLDN2\,
datab => \GRLFPC2_0.R.MK.RST_RET_6\,
datac => \GRLFPC2_0.R.MK.RST2\,
datad => \GRLFPC2_0.COMB.V.MK.RST_1_0_A2_3\);
GRLFPC2_0_COMB_UN3_IUEXEC: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC2_0.COMB.UN3_IUEXEC\,
dataa => \GRLFPC2_0.R.M.FPOP\,
datab => \GRLFPC2_0.R.X.FPOP\,
datac => \GRLFPC2_0.COMB.UN3_IUEXEC_0\);
GRLFPC2_0_R_A_FPOP_RNINLPU: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000000000000")
port map (
combout => \GRLFPC2_0.ANNULRES_0_SQMUXA_10\,
dataa => N_161,
datab => N_160,
datac => \GRLFPC2_0.R.A.FPOP\,
datad => \GRLFPC2_0.ANNULRES_0_SQMUXA_10_0\);
GRLFPC2_0_R_MK_BUSY2_RET_1_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.R.MK.BUSY2_RET_1_0_0_A2_0_G0\,
dataa => N_8,
datab => \GRLFPC2_0.R.MK.BUSY_RET_3\,
datac => \GRLFPC2_0.R.MK.BUSY_RET_4\,
datad => \GRLFPC2_0.COMB.V.MK.BUSY_2_4\);
GRLFPC2_0_COMB_LOCK_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => CPO_LDLOCKZ,
dataa => N_91,
datab => \GRLFPC2_0.R.STATE\(0),
datac => \GRLFPC2_0.R.STATE\(1),
datad => \GRLFPC2_0.COMB.LOCK_1_1_X\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_27_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_27\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_3_1\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_3_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84),
datab => N_34381_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A7_4_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_4\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A15_1\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_17_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_17\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => N_28709_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_1_1\(62),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O21\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_13_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_13\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => N_34381_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_13_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_12_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_12\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_2\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_7_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_7\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A25_1\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_13_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_6_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_6\(32),
dataa => N_28709_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_1_1\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O2\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A20_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A20\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O20_6\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O13_0\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O6_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011001010110010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O6\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_0_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_0\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_6_1\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_2\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_5_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_1_0\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_7_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_7\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8577_I_0_A2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0_0_A2_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_0_0_A2\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_3_1\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_2_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_2\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_1\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_4_1\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_0_0_A2_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_0_A2\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_12_0_A2\(62));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_3_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_1_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_2_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_2\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\(58),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_O2\(25));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_1_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_1\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_7_1\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_1_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_I_X2\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_4_2\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_1_0_A2_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_1_0_A2\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_4_1\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11846_I_I_I_X2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_12_0_A2\(62));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A14_6_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_6\(62),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_2\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O21\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A14_7_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_7\(62),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => N_33227_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_6_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_6\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_6_1\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_12_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_7_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_7\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_13_1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_11_2\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_10_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_10\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_13_1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_12_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_11_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_11\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_4_1\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_1_1\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_12_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_13_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_13\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_13_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_10_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_1\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_3_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_3\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_M2\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_5_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_5\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_14_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_1\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_10_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_10\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_14_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O2\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_0_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_0\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_16_2\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_8_1\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_M29\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_2_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_2\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_M2\(19),
datad => N_32980_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_4_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_4\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_16_1\(27),
datac => N_28871_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O13_0\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_7_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_7\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A26_1\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_8_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_8\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_8_1\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_1_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O13_0\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_9_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_9\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_16_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_16\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A15_1\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_21_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_21\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_1\(61),
datad => N_34072_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_24_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_24\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_1_1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_13_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_4_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_4\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_5_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_5\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A17_1\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_6_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_6\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83),
datab => N_33495_1,
datac => N_33157_1,
datad => N_28871_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_8_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_8\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A17_1\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_7_1\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_7_1\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A25_1\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_11_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_11\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_1\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_15_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_15\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_0\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_23_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_23\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_10_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8577_I_0_A2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_24_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_24\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => N_33157_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_2\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_25_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_25\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A17_1\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_7_1\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_2_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_2\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_7_1\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_M23\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_12_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_4_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_4\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_2\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_I_X2\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_6_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_6\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A22_1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_1\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_7_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_7_1\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_8_1\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0_1\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_8_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_8\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_7_1\(0),
datab => N_33157_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A25_1\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_10_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_10\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_1\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_12_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_11_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_10_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_12_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_16_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_16\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_8_1\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_12_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_18_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_18\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_16_1\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_7_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_20_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_20\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_2\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_3_1\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_O28_5\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0_1\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A28_3_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_3\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_13_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_12_1\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A28_9_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_9\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_3_1\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_2\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A28_11_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_11\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A28_15_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_15\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_2\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_1_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A28_16_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_16\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\(58),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A28_17_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_17\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A28_19_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_19\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_13_1\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A28_22_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_22\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_1\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_2\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_3_1\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A28_24_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_24\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_O28_5\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0_1\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_4_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_4\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_M26\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_12_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_5_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_5\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_1_1\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_7_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_7\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_6_1\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_8_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_8\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_2\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A25_1\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_9_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_9\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O18_4\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_11_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_11\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_1\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_5_1\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_12_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_12\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_0\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8577_I_0_A2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_21_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_21\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_1\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_11_2\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_22_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_22\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_M22\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_28_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_28\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_4_2\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_12_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_30_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_30\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_1_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_36_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_36\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_2\(25),
datac => N_33157_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_38_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_38\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_14_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_2\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O22_0_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110100011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_0\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_5_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_5\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_1_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_6_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_6\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_16_1\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O13_0\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_2_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_2\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_1_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_1\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_1\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_4_1\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_12_1\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_2_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000011000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_2\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_9_1\(0),
datac => N_29496_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_5_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_7_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_7\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_4_1\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_11_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_11\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78),
datab => N_33157_1,
datac => N_29496_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_12_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_12\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A17_1\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_14_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_14\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_0_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_0\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_1_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_M2_0\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_4_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_4\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_5_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_6_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001110100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_6\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_6_0\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_9_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_9\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_1_1\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_4_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_2\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_11_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_11\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A15_1\(18),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_1\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O25\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_16_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_16\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_16_1\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_9_1\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_2\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_19_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_19\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O25\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_20_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_20\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A19_1\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_7_1\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O2\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_2_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_2\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_M2_0\(6),
datad => N_34072_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_6_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_6\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O18_4\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(4),
datad => N_34072_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_8_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_8\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_10_1\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_14_1\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_9_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_9\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_10_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_4_1\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A26_1\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_10_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_10\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_2\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A24_1_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_1\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_M24\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A24_3_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_3\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_16_1\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A24_4_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_4\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN1_S_DYADIC_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A24_6_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_6\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_15_2\(60),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A24_13_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_13\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_3_1\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_1_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010100000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_1\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_M2\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_2\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_9_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_9\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_1\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_9_1\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_5_1\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_10_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_10\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_1_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_2\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_11_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_1_1\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_5_1\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_12_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_12\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_9_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O2\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_15_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_15\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O18_0\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_16_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_16\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O18_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O2\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_17_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_17\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_5_1\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_19_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_19\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_2_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000110100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_2\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80),
datab => N_28709_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_1\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_12_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_4_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_4\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0_1\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_5_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_5\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_8_1\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_1_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_3\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_8_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_8\(54),
dataa => N_28709_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_6_1\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0_1\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_9_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_9\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_16_2\(61),
datab => N_28709_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_11_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_11\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_2\(57),
datab => N_33157_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A25_1\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_13_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_13\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_16_2\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0_1\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_16_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_16\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_4_2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0_1\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_19_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_19\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80),
datac => N_33157_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0_1\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_21_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_21\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A17_1\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_23_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_23\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_2\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_24_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_24\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A7_1\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A17_1\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A26_1\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_4_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_4\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_4_2\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_5_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_5\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_2_1\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A26_1\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_6_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_6\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_7_1\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_2\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_1\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_6_1\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_8_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_8\(13),
dataa => N_33495_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_4_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_2\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_13_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_13\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_1_1\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_5_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_14_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_14\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A17_1\(34),
datab => N_32980_1,
datac => N_34072_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O2\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_15_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_15\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A17_1\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_1_1\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8577_I_0_A2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A30_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_1_1\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_8_1\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_12_1\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A30_2_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_2\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_1_1\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_12_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O25\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A30_3_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_3\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_13_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_1_1\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_7_1\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O13_0\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A30_4_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_4\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
datac => N_28709_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_5_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A30_6_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_6\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_1_1\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_8_1\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_14_1\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A30_7_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_7\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A22_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_13_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O2\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_16_1\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A30_8_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_8\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_5_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A30_11_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_11\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A30_13_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_13\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_8_1\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A30_16_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_16\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_1_1\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A30_17_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_17\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A30_18_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_18\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_14_1\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A30_22_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_22\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O13_0\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_2_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_2\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_7_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_5_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_8_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_8\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_8_0\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_1\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_9_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_9\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_14_1\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O13_0\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_10_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_10\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_14_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_2\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_15_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_15\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN1_S_DYADIC_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_4_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_4\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_M2\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_6_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_6\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84),
datab => N_33495_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_8_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_8\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(61),
datad => N_28871_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_9_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_9\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_2\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_16_1\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O21\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_10_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_10\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_2\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8577_I_0_A2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_11_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_11\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_16_1\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_1\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_12_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_12\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A3\(3),
datab => N_33157_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_12_1\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_15_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_15\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_16_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_16\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(13),
datad => N_28871_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_17_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_17\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_19_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_19\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_16_1\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_7_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_I_A26_2_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_2\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A3\(3),
datab => N_33157_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_16_1\(54),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O13_0\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_I_A26_7_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_7\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_I_A26_8_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_8\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O13_0\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_I_A26_9_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_9\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_2\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_16_1\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_I_A26_10_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_10\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_0\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_16_1\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_I_A26_12_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_12\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_13_1\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_I_X2\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_I_A26_13_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_13\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_10_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_2\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_I_X2\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_I_A26_14_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_14\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A13_1\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_I_A26_18_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_18\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_10_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_8_1\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_I_A26_19_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_19\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A28_1\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O13_0\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_I_A26_22_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_22\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O18_4\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\(19),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_16_1\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_I_A26_23_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_23\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O18_4\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_2\(57),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_12_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_1_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_1\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_1_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_4_1\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_14_1\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_7_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_7\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_13_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_14_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_14\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_9_1\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_3_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_3\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_3\(51),
datad => N_34072_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_4_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_2\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_1\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_5_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_5\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_7_1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O21\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_7_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_7\(51),
dataa => N_33227_2,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A15_1\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_1_1\(62),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O21\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_9_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_9\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A15_1\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O2\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_13_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_13_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_13\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_1_1\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O2\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_13_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_14_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_14\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_4_2\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A15_1\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A22_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O21\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_16_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_16\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_16_1\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_1_1\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_5_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_18_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_18\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A15_1\(18),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A22_1\(6),
datac => N_28871_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O2\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_1_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_1\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_M17\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_2_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_2\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84),
datab => N_33157_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_0\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_6_1\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_4_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_4\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_2\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN1_S_DYADIC_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_5_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_5\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => N_33157_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A7_3_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_3\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X3\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\(58),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O13_0\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_M2\(5),
datad => N_34072_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_2_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_2\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_M16\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_14_2\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_2_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_4_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_4\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_2\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_1_1\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_4_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_9_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_9\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_1_1\(62),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_0_2\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_10_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_10\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_16_1\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_10_0\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_12_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_12\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_16_1\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_1_1\(62),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_12_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_4_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_4\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_14_1\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_6_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_6\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O2\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_I_A26_5_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_5\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_1_1\(0),
datad => N_29496_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_I_A26_0_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_0\(31),
dataa => N_32980_1,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_2_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_3_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_3\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_10_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_1\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_1\(49),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_13_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A24_0_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_0\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_10_1\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_2\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_4_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_5_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_5\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_2\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_7_1\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_5_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_1_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_1\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_1_1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_3\,
datad => N_34072_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_23_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_23\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_2\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A28_2_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_2\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_13_1\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_2\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_1_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_1\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN1_S_DYADIC_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A25_1\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A29_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_16_1\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_2_A2_1_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_2_A2_1\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_14_1\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_1_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_1\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_2\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_5_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_5\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_9_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A19_1\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A25_1\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_2\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_4_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_4\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_10_1\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_14_1\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_4_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_4\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_0_I_O2\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_17_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_17\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_2\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_1_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_1\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datab => N_34381_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_0\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_14_1\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_46__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_2\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN1_S_DYADIC_0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_76_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_76__G0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(72),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN10_S_MOV: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN10_S_MOV\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_7_1\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_7_1\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_14_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_14\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_14_1\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O2\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_10_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_10\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_10_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O18_0\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_7_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_7\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A22_1\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_4_1\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_7_1\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_2\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_6_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_6\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A25_1\(27),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_8_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_8\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_9_1\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_1_1\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_14_1\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_17_1_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_17_1\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80),
datad => N_32980_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_7_1_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_7_1\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_1_3_TZ_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110111001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_3_TZ\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_12_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101010010010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2_2_TZ\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_13_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_13_1\(4));
GRLFPC2_0_V_FSR_AEXC_1_SQMUXA_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111100000000")
port map (
combout => \GRLFPC2_0.V.FSR.AEXC_1_SQMUXA_0\,
dataa => N_404,
datab => N_403,
datac => N_402,
datad => \GRLFPC2_0.V.FSR.NONSTD_0_SQMUXA_6_X\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_7_1\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_12_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_12\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_5_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_37_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_37\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datab => N_33227_2,
datac => N_29496_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_12_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_18_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_18\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83),
datac => N_33227_2,
datad => N_29496_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_0_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_1_0_0_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_1_0_0\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_2\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_4_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001001010010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2_5_TZ\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_1_TZ_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101010111011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_1_TZ\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_M27_0\(47),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_6_1\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_7_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001110001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2_5_TZ\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_3_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000001001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2_2_TZ\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_10_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2_9023_TZ\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_14_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000011000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2_8692_TZ\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011010011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011010011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN4_NOTAINFNAN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN4_NOTAINFNAN\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.EXPYBUS\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(239),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.EXPYBUS\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(238),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110101001101010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.EXPYBUS_0\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_V_0_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001110010010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011010011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(232),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_UN11_INFORCREGSN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLCREGXZ.UN11_INFORCREGSN\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.SELECTQUOBITS.NOTDIVC\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD57\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(1));
GRLFPC2_0_WRADDR_1_SQMUXA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101010100010101")
port map (
combout => \GRLFPC2_0.WRADDR_1_SQMUXA\,
dataa => \GRLFPC2_0.WRADDR_0_SQMUXA_X\,
datab => \GRLFPC2_0.R.I.V\,
datac => \GRLFPC2_0.R.X.FPOP\,
datad => \GRLFPC2_0.R.I.EXEC\);
GRLFPC2_0_COMB_V_I_EXEC_4_IV_0_A2_X_RNI5O6J1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111100000000")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.CEXC_1_SN_M2\,
dataa => N_404,
datab => N_403,
datac => N_402,
datad => \GRLFPC2_0.N_1570_I_I_A2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_114_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(114),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(117),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.ROMXZSL2FROMC\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(62),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(62));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(63),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(63),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(63));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_64_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(64),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(64),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(64));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_65_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(65),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(65));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_66_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(66),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(66),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(66));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_67_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(67),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(67),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(67));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_68_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(68),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(68),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(68));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_69_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(69),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(69),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(69));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_71_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(71),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(71),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(71));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_72_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(72),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(72),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(72));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_73_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(73),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(73),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(73));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_74_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(74),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(74),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(74));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(75),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(75),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(75));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_76_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(76),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(76),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(76));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_77_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(77),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(77),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(77));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_78_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_79_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_80_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_81_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_82_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(82));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_83_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_87_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(87),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(87),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(87));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_88_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(88),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(88),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(88));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_89_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(89),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(89),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(89));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_90_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(90),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(90),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(90));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_91_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(91),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(91),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(91));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_92_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(92),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(92),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(92));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_93_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(93),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(93),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(93));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_94_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(94),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(94),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(94));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_95_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(95),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(95),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(95));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_96_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(96),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(96),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(96));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_97_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(97),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(97),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(97));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_99_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(99),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(99),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(99));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_100_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(100),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(100),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(100));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_101_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(101),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(101),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(101));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_102_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(102),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(102),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(102));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_103_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(103),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(103),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(103));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_104_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(104),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(104),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(104));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_105_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(105),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(105),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(105));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_106_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(106),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(106),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(106));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_109_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(109),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(109),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(109));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_110_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(110),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(110),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(110));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_111_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(111),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(111),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(111));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_112_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(112),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(112),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(112));
\GRLFPC2_0_WRDATA_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(10),
dataa => N_402,
datab => N_420,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(42));
\GRLFPC2_0_WRDATA_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(3),
dataa => N_402,
datab => N_413,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(35));
\GRLFPC2_0_WRDATA_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(2),
dataa => N_402,
datab => N_412,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(34));
\GRLFPC2_0_WRDATA_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(10),
dataa => N_402,
datab => N_420,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(10));
\GRLFPC2_0_WRDATA_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(3),
dataa => N_402,
datab => N_413,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(3));
\GRLFPC2_0_WRDATA_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(2),
dataa => N_402,
datab => N_412,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(2));
\GRLFPC2_0_WRDATA_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(0),
dataa => N_402,
datab => N_410,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(0));
\GRLFPC2_0_WRDATA_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(28),
dataa => N_402,
datab => N_438,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(60));
\GRLFPC2_0_WRDATA_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(7),
dataa => N_402,
datab => N_417,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(39));
\GRLFPC2_0_WRDATA_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(9),
dataa => N_402,
datab => N_419,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(9));
\GRLFPC2_0_WRDATA_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(7),
dataa => N_402,
datab => N_417,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(7));
\GRLFPC2_0_WRDATA_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(19),
dataa => N_402,
datab => N_429,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(51));
\GRLFPC2_0_WRDATA_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(16),
dataa => N_402,
datab => N_426,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(48));
\GRLFPC2_0_WRDATA_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(13),
dataa => N_402,
datab => N_423,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(45));
\GRLFPC2_0_WRDATA_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(28),
dataa => N_402,
datab => N_438,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(28));
\GRLFPC2_0_WRDATA_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(19),
dataa => N_402,
datab => N_429,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(19));
\GRLFPC2_0_WRDATA_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(16),
dataa => N_402,
datab => N_426,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(16));
\GRLFPC2_0_WRDATA_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(13),
dataa => N_402,
datab => N_423,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(13));
\GRLFPC2_0_WRDATA_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011110000")
port map (
combout => RFI1_WRDATAZ(31),
dataa => N_402,
datab => N_441,
datac => \GRLFPC2_0.WRDATA_0_X\(63),
datad => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\);
\GRLFPC2_0_WRDATA_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(23),
dataa => N_402,
datab => N_433,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(55));
\GRLFPC2_0_WRDATA_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(20),
dataa => N_402,
datab => N_430,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(52));
\GRLFPC2_0_WRDATA_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(17),
dataa => N_402,
datab => N_427,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(49));
\GRLFPC2_0_WRDATA_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(14),
dataa => N_402,
datab => N_424,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(46));
\GRLFPC2_0_WRDATA_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(11),
dataa => N_402,
datab => N_421,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(43));
\GRLFPC2_0_WRDATA_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(8),
dataa => N_402,
datab => N_418,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(40));
\GRLFPC2_0_WRDATA_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(31),
dataa => N_402,
datab => N_441,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(31));
\GRLFPC2_0_WRDATA_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(23),
dataa => N_402,
datab => N_433,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(23));
\GRLFPC2_0_WRDATA_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(20),
dataa => N_402,
datab => N_430,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(20));
\GRLFPC2_0_WRDATA_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(17),
dataa => N_402,
datab => N_427,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(17));
\GRLFPC2_0_WRDATA_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(14),
dataa => N_402,
datab => N_424,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(14));
\GRLFPC2_0_WRDATA_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(11),
dataa => N_402,
datab => N_421,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(11));
\GRLFPC2_0_WRDATA_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(8),
dataa => N_402,
datab => N_418,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(8));
\GRLFPC2_0_WRDATA_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(30),
dataa => N_402,
datab => N_440,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(62));
\GRLFPC2_0_WRDATA_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(27),
dataa => N_402,
datab => N_437,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(59));
\GRLFPC2_0_WRDATA_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(25),
dataa => N_402,
datab => N_435,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(57));
\GRLFPC2_0_WRDATA_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(30),
dataa => N_402,
datab => N_440,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(30));
\GRLFPC2_0_WRDATA_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(27),
dataa => N_402,
datab => N_437,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(27));
\GRLFPC2_0_WRDATA_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(25),
dataa => N_402,
datab => N_435,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(25));
\GRLFPC2_0_WRDATA_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(6),
dataa => N_402,
datab => N_416,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(38));
\GRLFPC2_0_WRDATA_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(5),
dataa => N_402,
datab => N_415,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(37));
\GRLFPC2_0_WRDATA_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(6),
dataa => N_402,
datab => N_416,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(6));
\GRLFPC2_0_WRDATA_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(5),
dataa => N_402,
datab => N_415,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(5));
\GRLFPC2_0_WRDATA_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(24),
dataa => N_402,
datab => N_434,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(56));
\GRLFPC2_0_WRDATA_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(12),
dataa => N_402,
datab => N_422,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(44));
\GRLFPC2_0_WRDATA_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(0),
dataa => N_402,
datab => N_410,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(32));
\GRLFPC2_0_WRDATA_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(24),
dataa => N_402,
datab => N_434,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(24));
\GRLFPC2_0_WRDATA_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(12),
dataa => N_402,
datab => N_422,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(12));
\GRLFPC2_0_WRADDR_1_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRADDRZ(3),
dataa => N_402,
datab => N_409,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.COMB.WRADDR_5_X\(4));
\GRLFPC2_0_WRDATA_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(21),
dataa => N_402,
datab => N_431,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(53));
\GRLFPC2_0_WRDATA_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(18),
dataa => N_402,
datab => N_428,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(50));
\GRLFPC2_0_WRDATA_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(15),
dataa => N_402,
datab => N_425,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(47));
\GRLFPC2_0_WRDATA_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(21),
dataa => N_402,
datab => N_431,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(21));
\GRLFPC2_0_WRDATA_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(18),
dataa => N_402,
datab => N_428,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(18));
\GRLFPC2_0_WRDATA_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(15),
dataa => N_402,
datab => N_425,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(15));
\GRLFPC2_0_WRDATA_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(1),
dataa => N_402,
datab => N_411,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(33));
\GRLFPC2_0_WRDATA_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(22),
dataa => N_402,
datab => N_432,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(22));
\GRLFPC2_0_WRDATA_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(1),
dataa => N_402,
datab => N_411,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(1));
\GRLFPC2_0_WRDATA_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(29),
dataa => N_402,
datab => N_439,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(61));
\GRLFPC2_0_WRDATA_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(4),
dataa => N_402,
datab => N_414,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(36));
\GRLFPC2_0_WRDATA_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(29),
dataa => N_402,
datab => N_439,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(29));
\GRLFPC2_0_WRDATA_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(4),
dataa => N_402,
datab => N_414,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(4));
\GRLFPC2_0_WRDATA_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(22),
dataa => N_402,
datab => N_432,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(54));
\GRLFPC2_0_WRADDR_1_I_M2_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRADDRZ(2),
dataa => N_402,
datab => N_408,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.COMB.WRADDR_5_I_M2_X\(3));
\GRLFPC2_0_WRADDR_1_I_M2_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRADDRZ(1),
dataa => N_402,
datab => N_407,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.COMB.WRADDR_5_I_M2_X\(2));
\GRLFPC2_0_WRADDR_1_I_M2_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRADDRZ(0),
dataa => N_402,
datab => N_406,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.COMB.WRADDR_5_I_M2_X\(1));
\GRLFPC2_0_WRDATA_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(26),
dataa => N_402,
datab => N_436,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(58));
\GRLFPC2_0_WRDATA_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI1_WRDATAZ(9),
dataa => N_402,
datab => N_419,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(41));
\GRLFPC2_0_WRDATA_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111110000000")
port map (
combout => RFI2_WRDATAZ(26),
dataa => N_402,
datab => N_436,
datac => \GRLFPC2_0.COMB.UN31_DEBUG_UNIT_X\,
datad => \GRLFPC2_0.WRDATA_0_X\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000101000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001101000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(133),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(17),
datac => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(122),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(6),
datac => \GRLFPC2_0.FPI.LDOP_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(119),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(3),
datac => \GRLFPC2_0.FPI.LDOP_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(20));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_A_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_A_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(120),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(4),
datac => \GRLFPC2_0.FPI.LDOP_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_A\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_A_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_A\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(121),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(5),
datac => \GRLFPC2_0.FPI.LDOP_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(129),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(13),
datac => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(132),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(16),
datac => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(130),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(14),
datac => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(141),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1_X\(25),
datac => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(140),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1_X\(24),
datac => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(128),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(12),
datac => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(126),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(10),
datac => \GRLFPC2_0.FPI.LDOP_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(134),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(18),
datac => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(21),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(137),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(21),
datac => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(25));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(138),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(22),
datac => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(139),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1_X\(23),
datac => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(123),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(7),
datac => \GRLFPC2_0.FPI.LDOP_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(127),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(11),
datac => \GRLFPC2_0.FPI.LDOP_REP2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN15_XZROUNDOUT\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(124),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(8),
datac => \GRLFPC2_0.FPI.LDOP_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(46),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(40),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(50));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(136),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(20),
datac => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_235_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000010101010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0\(235),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.FPI.OP2_X\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPAREGLOADEN\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(16),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011101000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.UN17_U_RDN\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(21),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_A\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_A_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111100110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_A\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_A_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(38));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(40),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(40));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(45),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_A_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(45),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_A_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(43),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(43),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(45),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(35));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(35));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_A_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_A_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(21),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(20),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(14));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(20),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010111100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_A\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_A_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001100101011101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12_A\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(25));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_A_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_A_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(21),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_A_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(21),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_A_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_A_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_A_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_A_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(35));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_A_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_A_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_A_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_A_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(22),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(28));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(40),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(131),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(15),
datac => \GRLFPC2_0.FPI.LDOP_REP2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(46),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS_2\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100011011000110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100011011000110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP2\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0_REP1\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100011011000110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100011011000110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116_REP1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0_REP1\(0));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0_REP1\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(46),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(35));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_A_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_A_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_3_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_2\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_3_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_2\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(16),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_3_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000011100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(255),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3_A\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_3_A_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3_A\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN8_TEMP_U_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN8_TEMP_U\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN8_TEMP_2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(50));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_A_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_A_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_A_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_A_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_A_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_0_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_0\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_0_A\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_0_A_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_0_A\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_0_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_0\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_0_A\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_0_A_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_0_A\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_12\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_0_0_2__G0\,
dataa => N_69,
datab => N_66,
datac => N_68,
datad => N_64);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_0_0_1__G0\,
dataa => N_69,
datab => N_66,
datac => N_68,
datad => N_64);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000011111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW_6_0_0__G0\,
dataa => N_65,
datab => N_69,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW_6_0_0__G2_0_X\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MAPMULXFF.UN4_UNIMPMAP_X\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_372_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100110001001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_372__G1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0_REP2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_2\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.SELINITREMBIT\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_GRFPUF_0_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF_0\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.SELINITREMBIT\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD52\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_GRFPUF_0_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF_0\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.SELINITREMBIT\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD53\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_GRFPUF_0_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF_0\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.SELINITREMBIT\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD54\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_GRFPUF_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011101000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.SELINITREMBIT\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD55\);
\GRLFPC2_0_R_I_CC_RNO_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000000010")
port map (
combout => \GRLFPC2_0.R.I.CC_0_0_1__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(39),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(40));
\GRLFPC2_0_R_I_CC_RNO_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100000")
port map (
combout => \GRLFPC2_0.R.I.CC_0_0_0__G2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(39),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(40));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXCEP_1_TZ_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000011100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.EXCEP_1_TZ\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(40),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(39));
GRLFPC2_0_COMB_FPDECODE_ST_0_A2_0_A2_0_X_RNI97AM: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.R.A.ST_RET_0_0_G1\,
dataa => N_87,
datab => N_80,
datac => N_88,
datad => \GRLFPC2_0.COMB.FPDECODE.ST_0_A2_0_A2_0_X\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_RNIGFVI_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010101000101010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6));
GRLFPC2_0_COMB_V_FSR_RD_1_SN_M2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111100000000")
port map (
combout => \GRLFPC2_0.COMB.V.FSR.RD_1_SN_M2\,
dataa => N_404,
datab => N_403,
datac => N_402,
datad => N_8);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNI0VD2_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000011100000")
port map (
combout => G_8368,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLOADEN_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLAREGEXP.EXPAREGLOADEN_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(47),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD12\,
datac => \GRLFPC2_0.FPI.LDOP_REP0\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_A_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_A\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP2\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111000001110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_108_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(108),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(108),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(108));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_107_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(107),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(107),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(107));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_98_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(98),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(98),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(98));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_86_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(86),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(86),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(86));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIB5V7_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101001011010010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN6_NOTPROP_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(371),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_RNII9BI_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111000001110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULLSBLOGIC.TEMP_2\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(50));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(43),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_0_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(45),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(125),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(9),
datac => \GRLFPC2_0.FPI.LDOP_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M3_70_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(70),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(70),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(70));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_UN4_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.UN4_TEMP2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(72),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(63));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CONDMUXMULXFF_UN4_NOTSQRTLFTCC: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CONDMUXMULXFF.UN4_NOTSQRTLFTCC\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(72),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIRP6Q_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G_32\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(51),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(49));
GRLFPC2_0_R_X_AFSR_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC2_0.R.X.AFSR_0_0_G1\,
dataa => N_299,
datab => N_298,
datac => \GRLFPC2_0.R.M.AFQ_RET_1\,
datad => \GRLFPC2_0.R.M.AFSR_RET\);
GRLFPC2_0_R_X_AFQ_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC2_0.R.X.AFQ_0_0_G1\,
dataa => N_299,
datab => N_298,
datac => \GRLFPC2_0.R.M.AFQ_RET_1\,
datad => \GRLFPC2_0.R.M.AFQ_RET\);
GRLFPC2_0_R_X_FPOP_RNIAQIJ: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC2_0.R.I.RDD_0_0_G1_0_8238_I_O4\,
dataa => N_368,
datab => N_367,
datac => N_18,
datad => \GRLFPC2_0.R.X.FPOP\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M13_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M11\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M8\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M11S4\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M13_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M11\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M8\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M11S4\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M12_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M2\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5S4\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M12_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M2\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5S4\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_0_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100000110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.EXPYBUS_0\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2_1\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100111001001110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(241),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2_1\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_0_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100000110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.EXPYBUS_0\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2_1\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_0_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100000110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.EXPYBUS_0\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(237),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2_1\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_236_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000010101010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0\(236),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datac => \GRLFPC2_0.FPI.OP2_X\(60),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPAREGLOADEN\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_1_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_1\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_115_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(115),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(118),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.ROMXZSL2FROMC\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(135),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(19),
datac => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_2_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_2\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_9_0_A2\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_3_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_3\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O2\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_1_0\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_RNISLCO3_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_9\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(48),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_27_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_27\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_18_2\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_7_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_7\(62),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_26_2\(60),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_9_0_A2\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_12_0_A2\(62),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_14_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_14\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_7_1\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_5_0_A2_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_5_0_A2\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_12_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_6_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_6\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_1_0\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_1_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_1\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_4_1\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0_A2_0_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_0_A2_0\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80),
datac => N_34381_1,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_O2\(25));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_7_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_7\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_14_2\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2\(40),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_26_2\(60),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_4_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_4\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN1_S_DYADIC_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_12_0_A2_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_12_0_A2\(62),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_9_0_A2_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_9_0_A2\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_0_A2_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_0_A2\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_8_0_A2_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_8_0_A2\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_30_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_30\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O18_4\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_22_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_22\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O18_4\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_0_A2_1_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_A2_1\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_14_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_14\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_8_1\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_3_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datab => N_34381_1,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(4),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_1_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_1\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_2\(25),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_4785_A2_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A28_11_0_A2_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_A28_11_0_A2\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_23_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_23\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_45_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_45\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_2_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111000111110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_2\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11_2\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O6_1_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111000100001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O6_1\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O6_2_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000110000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O6_2\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O20_5_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000011000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O20_5\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O7_0_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100110000011101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O7_0\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O7_1_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001100001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O7_1\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O7_2_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010001110001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O7_2\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_O16_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000110100001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O16\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O16_1_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101100001011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_1\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O23_7_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101100001011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_7\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O23_8_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001110000011100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_8\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O23_8_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_8\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_O28_6_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110110101101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_O28_6\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_0_M2_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110000111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_M2\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O26_8_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010010100100101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O26_8\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O26_9_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001000110010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O26_9\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O22_11_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000000100011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_11\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_O27_4_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011100100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_O27_4\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_O24_3_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_O24_3\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O23_6_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110010001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_6\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O19_4_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100001001000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_4\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_O13_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100001001000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_O13\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O17_1_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010000110100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O17_1\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O16_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000110000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_10_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_10\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_2_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_2\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_4\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_13_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_13\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_21_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_21\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O18_0\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A28_14_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_14\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_5_1\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_2_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_2\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_2_3\(18),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_16_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_16\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_14_2\(59),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_5_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_5\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83),
datad => N_34072_1);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_11_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_11\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_4_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_13_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_13\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(13),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_13_1\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_16_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_16\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_2\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_5_1\(6),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_14_1\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_22_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_22\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_16_1\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O21\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_I_A26_16_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_16\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_6_1\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_10_2_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_10_2\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A15_1\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_5_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_5\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_0\(5),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_5_1\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_14_0_A2_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_14_0_A2\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_26_2\(60));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_1_A2_1_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1_A2_1\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_1_0_A2\(62));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_11_0_A2_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_11_0_A2\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_4_2\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_4_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_4\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_12_0_A2\(62));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_7_1\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN1_S_DYADIC_0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(61),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIN7RL_71_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011111101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(72),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(71),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_2_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010011000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_2_SQMUXA_2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLBREGXZ.UN4_XZBREGLOADEN\,
datac => \GRLFPC2_0.FPI.LDOP_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CHECKOVANDDENORM_UN13_NOTPOSSIBLEOV_4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD49\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD50\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD54\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CHECKOVANDDENORM_UN13_NOTPOSSIBLEOV_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD47\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD48\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD53\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN30_CONDITIONAL_M2_E_4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN30_CONDITIONAL_M2_E_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD3\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD5\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD6\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN30_CONDITIONAL_M2_E_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN30_CONDITIONAL_M2_E_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD7\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN10_U_SNNOTDB_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.UN10_U_SNNOTDB_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(10),
datac => \GRLFPC2_0.FPI.LDOP_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN17_SHDVAR_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A7_0_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A7_0\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_2_0_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_2_0\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A22_0_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A22_0\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIJ3LJ_73_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101000011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.TEMP_25_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(74),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(72),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_2_0_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100110001001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_2_0\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_12_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2_8645_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_3_1_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001100000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_1\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_7_0_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_7_0\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_6_0_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_6_0\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_3_1_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_3_1\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_9_0_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010101000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_9_0\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_0_0_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_0_0\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_13_0_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_13_0\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_0_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0_0\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A24_7_0_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_7_0\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_1_1_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101110001011100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_1_1\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_5_0_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_5_0\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_8_0_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010000010100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_8_0\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_2_0_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_2_0\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A25_1\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A14_2_2_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011101100111011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_2_2\(62),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_3_1_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011101000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_3_1\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_11_0_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000010110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11_0\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A30_1_0_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_1_0\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_23_0_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_23_0\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A24_11_0_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_11_0\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A24_5_0_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_5_0\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A28_23_0_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_23_0\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_12_0_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_12_0\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN12_SRTOSTICKY_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN12_SRTOSTICKY_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD6\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD7\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD8\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD9\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_5_0_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_5_0\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_7_0_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000101000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7_0\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_5_0_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_5_0\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_11_0_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_11_0\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_10_1_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_10_1\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_15_0_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_15_0\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_4_0_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_4_0\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_2_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0_2\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_6_0_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_6_0\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_0_0_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0_0\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_2_0_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_2_0\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_1_0_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_1_0\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_9_0_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_9_0\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_10_1_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_10_1\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83));
GRLFPC2_0_COMB_V_A_AFSR_1_1_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC2_0.COMB.V.A.AFSR_1_1_0\,
dataa => \GRLFPC2_0.R.A.AFQ_RET\(7),
datab => \GRLFPC2_0.R.A.MOV_RET\(12),
datac => \GRLFPC2_0.R.A.MOV_RET\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_15_0_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_15_0\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_0_11_0_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0_11_0\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_10_0_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_10_0\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O29_1_0_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010100010101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O29_1_0\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A28_25_1_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_25_1\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A28_25_0_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_25_0\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_5_0_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_5_0\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_2_0_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_2_0\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_10_1_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_10_1\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN3_S_SQRT_1_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_1_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_0_0_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_0_0\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_16_1_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_16_1\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_16_0_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_16_0\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_5_0_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_5_0\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_3_0_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_3_0\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_5_0_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_0\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_17_1_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000110100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_17_1\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_17_0_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_17_0\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_12_0_0_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_12_0_0\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_16_0_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_16_0\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_10_0_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_10_0\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_3_1_0_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_3_1_0\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_17_1_0_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_17_1_0\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_6_1_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000010100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_6_1\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_20_0_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_20_0\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A30_10_0_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000010100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_10_0\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A7_4_0_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_4_0\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_I_A26_4_0_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_4_0\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A28_1\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A24_9_1_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_9_1\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A24_9_0_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_9_0\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_3_1_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_3_1\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_3_0_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_3_0\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_18_1_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_18_1\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_20_0_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_20_0\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_11_1_0_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_11_1_0\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_11_0_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_11_0\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A30_21_0_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_21_0\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A14_0_1_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_0_1\(62),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A14_0_0_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_0_0\(62),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_22_1_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_22_1\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A30_27_1_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_27_1\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_4_0_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001100000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_4_0\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_14_0_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101000011010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_14_0\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_12_0_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110000001100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_12_0\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_11_0_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011000000110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_11_0\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_I_A26_21_1_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_21_1\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_13_1_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_13_1\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A30_5_0_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_5_0\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_12_0_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_12_0\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_20: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_20\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_19: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_19\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_17: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_17\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_16: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_16\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_15: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_15\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_14: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_14\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_I_A26_20_1_0_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_20_1_0\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_19_0_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_19_0\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_10_0_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_10_0\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_8_0_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_8_0\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_2_1_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_2_1\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_O2_1_0_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011001000110010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_O2_1_0\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A28_6_0_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A28_6_0\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_3_0_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000010010000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_3_0\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_6_0_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_6_0\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83));
GRLFPC2_0_R_A_LD_RNI5CHL: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.COMB.FPOP_0_0_O2_0_2\,
dataa => \GRLFPC2_0.R.A.LD\,
datab => \GRLFPC2_0.R.E.LD\,
datac => \GRLFPC2_0.R.M.LD\,
datad => \GRLFPC2_0.R.X.LD\);
GRLFPC2_0_COMB_UN1_MEXC_1_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011101110111")
port map (
combout => \GRLFPC2_0.COMB.UN1_MEXC_1_1\,
dataa => \GRLFPC2_0.R.FSR.TEM\(1),
datab => \GRLFPC2_0.R.I.EXC\(1),
datac => \GRLFPC2_0.R.FSR.TEM\(0),
datad => \GRLFPC2_0.R.I.EXC\(0));
GRLFPC2_0_COMB_UN1_MEXC_1_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011101110111")
port map (
combout => \GRLFPC2_0.COMB.UN1_MEXC_1_0\,
dataa => \GRLFPC2_0.R.FSR.TEM\(3),
datab => \GRLFPC2_0.R.I.EXC\(3),
datac => \GRLFPC2_0.R.FSR.TEM\(2),
datad => \GRLFPC2_0.R.I.EXC\(2));
GRLFPC2_0_COMB_V_A_AFQ_1_7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.COMB.V.A.AFQ_1_7\,
dataa => \GRLFPC2_0.R.A.MOV_RET\(12),
datab => \GRLFPC2_0.R.A.AFQ_RET\(7),
datac => \GRLFPC2_0.R.A.MOV_RET\(13),
datad => \GRLFPC2_0.R.A.MOV_RET\(0));
GRLFPC2_0_COMB_V_A_AFQ_1_6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC2_0.COMB.V.A.AFQ_1_6\,
dataa => \GRLFPC2_0.R.A.MOV_RET\(11),
datab => \GRLFPC2_0.R.A.MOV_RET\(15),
datac => \GRLFPC2_0.R.A.AFQ_RET_2\,
datad => \GRLFPC2_0.R.A.AFQ_RET\(5));
GRLFPC2_0_COMB_V_MK_RST_1_0_A2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.COMB.V.MK.RST_1_0_A2_3\,
dataa => \GRLFPC2_0.R.MK.RST_RET_3\,
datab => \GRLFPC2_0.R.MK.RST_RET_2\,
datac => \GRLFPC2_0.R.MK.RST_RET\,
datad => \GRLFPC2_0.R.MK.LDOP_RET\);
GRLFPC2_0_COMB_UN2_HOLDN_0_A2_13_4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_13_4\,
dataa => \GRLFPC2_0.R.A.MOV_RET\(2),
datab => \GRLFPC2_0.R.A.MOV_RET\(10),
datac => \GRLFPC2_0.R.A.MOV_RET\(3),
datad => \GRLFPC2_0.R.A.MOV_RET\(8));
GRLFPC2_0_COMB_UN2_HOLDN_0_A2_13_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_13_3\,
dataa => \GRLFPC2_0.R.A.AFQ_RET\(9),
datab => \GRLFPC2_0.R.A.MOV_RET\(7),
datac => \GRLFPC2_0.R.A.MOV_RET\(6));
GRLFPC2_0_R_E_SEQERR_RNO_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.COMB.SEQERR.UN3_QNE_2\,
dataa => \GRLFPC2_0.R.A.AFQ_RET\(7),
datab => \GRLFPC2_0.R.A.MOV_RET\(11),
datac => \GRLFPC2_0.R.A.MOV_RET\(0),
datad => \GRLFPC2_0.R.A.AFQ_RET\(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN26_NOTAINFNAN_5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN26_NOTAINFNAN_5\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(237),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN26_NOTAINFNAN_4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN26_NOTAINFNAN_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(238),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(239),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(240),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(241));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN26_NOTBINFNAN_5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN26_NOTBINFNAN_5\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(250),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(257),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(255),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(256));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN26_NOTBINFNAN_4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN26_NOTBINFNAN_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(251),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(252),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(253),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(254));
GRLFPC2_0_N_939_I_I_A2_0_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100010")
port map (
combout => \GRLFPC2_0.N_939_I_I_A2_0_0\,
dataa => N_87,
datab => N_80,
datac => N_76,
datad => N_77);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN38_SHDVAR_3_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_3_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN38_SHDVAR_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55));
GRLFPC2_0_RIN_MK_LDOP_8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC2_0.RIN.MK.LDOP_8\,
dataa => \GRLFPC2_0.R.MK.LDOP_RET_1\(2),
datab => \GRLFPC2_0.R.MK.LDOP_RET_1\(6),
datac => \GRLFPC2_0.R.MK.LDOP_RET_1\(4),
datad => \GRLFPC2_0.R.MK.LDOP_RET\);
GRLFPC2_0_RIN_MK_LDOP_7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC2_0.RIN.MK.LDOP_7\,
dataa => \GRLFPC2_0.R.MK.LDOP_RET_1\(8),
datab => \GRLFPC2_0.R.MK.LDOP_RET_1\(7),
datac => \GRLFPC2_0.R.MK.LDOP_RET_1\(5),
datad => \GRLFPC2_0.R.MK.LDOP_RET_1\(1));
GRLFPC2_0_RIN_MK_LDOP_6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100000001")
port map (
combout => \GRLFPC2_0.RIN.MK.LDOP_6\,
dataa => \GRLFPC2_0.R.MK.LDOP_RET_3\,
datab => \GRLFPC2_0.R.MK.LDOP_RET_6\,
datac => \GRLFPC2_0.R.MK.LDOP_RET_4\(0),
datad => \GRLFPC2_0.R.MK.LDOP_RET_4\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNI9E7I_237_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_5\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(237),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNI8A7I_238_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_4\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(238),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(239),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(240),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(241));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIQ28I_250_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_5\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(250),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(257),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(255),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(256));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNII28I_251_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_4\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(251),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(252),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(253),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(254));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN9_WQSTSETS_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111011111110111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN9_WQSTSETS_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD4\);
GRLFPC2_0_V_FSR_FTT_1_SQMUXA_3_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000110100001101")
port map (
combout => \GRLFPC2_0.V.FSR.FTT_1_SQMUXA_3_0\,
dataa => \GRLFPC2_0.R.X.AFSR\,
datab => \GRLFPC2_0.R.X.LD\,
datac => \GRLFPC2_0.R.X.SEQERR\);
GRLFPC2_0_R_MK_BUSY_RET_4_RNO_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.R.MK.BUSY_RET_4_0_0_A2_0_G0_2\,
dataa => \GRLFPC2_0.R.MK.RST_RET_6\,
datab => \GRLFPC2_0.R.MK.RST2\,
datac => \GRLFPC2_0.R.MK.RST_RET\,
datad => \GRLFPC2_0.R.MK.LDOP_RET\);
GRLFPC2_0_COMB_UN4_LOCK_0_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC2_0.COMB.UN4_LOCK_0_2\,
dataa => \GRLFPC2_0.R.A.AFQ_RET_2\,
datab => \GRLFPC2_0.R.A.ST_RET_2\(1),
datac => \GRLFPC2_0.R.A.AFQ_RET_5\,
datad => \GRLFPC2_0.R.A.ST_RET_2\(0));
GRLFPC2_0_RS2_0_SQMUXA_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.RS2_0_SQMUXA_2\,
dataa => \GRLFPC2_0.R.A.AFQ_RET\(9),
datab => \GRLFPC2_0.R.A.MOV_RET\(12),
datac => \GRLFPC2_0.R.A.MOV_RET\(13),
datad => \GRLFPC2_0.R.A.MOV_RET\(15));
GRLFPC2_0_COMB_UN3_IUEXEC_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC2_0.COMB.UN3_IUEXEC_0\,
dataa => \GRLFPC2_0.R.E.FPOP\,
datab => \GRLFPC2_0.R.I.EXEC\,
datac => \GRLFPC2_0.R.A.FPOP\);
GRLFPC2_0_R_E_FPOP_RNI9JVD: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC2_0.ANNULRES_0_SQMUXA_10_0\,
dataa => \GRLFPC2_0.R.M.FPOP\,
datab => \GRLFPC2_0.R.X.FPOP\,
datac => \GRLFPC2_0.R.E.FPOP\,
datad => \GRLFPC2_0.R.I.EXEC\);
GRLFPC2_0_COMB_UN8_CCV_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010001000")
port map (
combout => \GRLFPC2_0.COMB.UN8_CCV_1\,
dataa => N_283,
datab => \GRLFPC2_0.R.M.FPOP\,
datac => \GRLFPC2_0.R.I.EXEC\,
datad => \GRLFPC2_0.R.I.INST\(19));
GRLFPC2_0_COMB_UN8_CCV_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010001000")
port map (
combout => \GRLFPC2_0.COMB.UN8_CCV_0\,
dataa => N_214,
datab => \GRLFPC2_0.R.E.FPOP\,
datac => \GRLFPC2_0.R.X.AFSR\,
datad => \GRLFPC2_0.R.X.LD\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_TOGGLESIG: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.TOGGLESIG\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(20),
datac => \GRLFPC2_0.FPI.LDOP_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN8_NOTBINFNAN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN8_NOTBINFNAN\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(249),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(247));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN3_NOTBZERODENORM: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN3_NOTBZERODENORM\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(249),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(247));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELINITREMBIT: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.SELINITREMBIT\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD56_RNI4E2D: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD54\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD55\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD56\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN17_U_RDN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.UN17_U_RDN\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(1),
datab => \GRLFPC2_0.R.FSR.RD\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(21),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_COMPUTECONST_UN25_RESVEC: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNI0V32_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.NOTAM2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.U_RDN_1_8221\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(2),
datab => \GRLFPC2_0.R.FSR.RD\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(21),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.UN17_U_RDN_I_0_8204_I_A2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(21),
datab => \GRLFPC2_0.R.FSR.RD\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(1));
GRLFPC2_0_RS2_0_SQMUXA_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC2_0.RS2_0_SQMUXA_3\,
dataa => \GRLFPC2_0.R.A.AFQ_RET\(7),
datab => \GRLFPC2_0.R.A.AFQ_RET\(5),
datac => \GRLFPC2_0.R.A.MOV_RET\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_173_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_68_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.WQSCTRL\(68),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(47),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD12\,
datac => \GRLFPC2_0.FPI.LDOP_REP5\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN4_NOTSHIFTCOUNT1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN4_NOTSHIFTCOUNT1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(14),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP2_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.TEMP2_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(72),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(71),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65));
GRLFPC2_0_COMB_V_MK_BUSY_2_4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.COMB.V.MK.BUSY_2_4\,
dataa => \GRLFPC2_0.R.MK.BUSY2_RET\,
datab => \GRLFPC2_0.R.MK.BUSY_RET_2\,
datac => \GRLFPC2_0.R.MK.BUSY_RET_5\,
datad => \GRLFPC2_0.R.MK.BUSY_RET\);
GRLFPC2_0_COMB_UN1_R_I_V_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001000")
port map (
combout => \GRLFPC2_0.COMB.UN1_R.I.V_0\,
dataa => \GRLFPC2_0.R.I.V\,
datab => \GRLFPC2_0.R.X.FPOP\,
datac => \GRLFPC2_0.R.I.EXEC\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN3_NOTAZERODENORM: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.AEBEEXC.UN3_NOTAZERODENORM\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234));
GRLFPC2_0_RS1D_CNST_0_A3_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.RS1D_CNST_0_A3_0\,
dataa => N_77,
datab => N_87,
datac => N_76,
datad => N_80);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_59__G0_YY\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
datab => \GRLFPC2_0.FPI.LDOP_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD54\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_1_0_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_1_0\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A15_0_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A15_0\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_0_0_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_0_0\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A13_0_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A13_0\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_17_0_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_17_0\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_7_0_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7_0\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_6_1_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_6_1\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_6_0_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_6_0\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_9_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_9_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_15_1_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_15_1\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_3_1_0_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_1_0\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_3_0_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_0\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A14_5_1_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_5_1\(62),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_8_1_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_8_1\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_14_0_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_14_0\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_9_0_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010101000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_9_0\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A14_1_1_0_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_1_1_0\(62),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_11_0_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_11_0\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_4_1_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_4_1\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_18_1_0_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_18_1_0\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_12_0_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_12_0\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_9_0_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_9_0\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83));
GRLFPC2_0_COMB_RDD_1_M14_0_A2_2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC2_0.COMB.RDD_1.M14_0_A2_2_1\,
dataa => N_65,
datab => N_64,
datac => N_66,
datad => N_76);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_22_0_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_22_0\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_7_0_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010100000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_7_0\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(314),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_3_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(247),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_3_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(260),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(258),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(263),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(262),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_4_0_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010111001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_4_0\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(311),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(289),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(282),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(298),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_TEMP: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100011111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SFTLFT.UN4_TEMP\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_TEMP: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110011101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(21),
datab => \GRLFPC2_0.FPI.LDOP_REP1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_3_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(232),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(245),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTDECODEDUNIMP_A_RNO_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN6_S\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(21),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(294),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(292),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(291),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(290),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(288),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(287),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(286),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(285),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(284),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(281),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_2_0_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011110111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_2_0\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(278),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(40),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(275),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110111111101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(259),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(295),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(279),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(293),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(264),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(266),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(304),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(274),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(273),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(45),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(270),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(268),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(306),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(301),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(297),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(300),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_UN129_TEMP_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011110111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.UN129_TEMP_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_UN126_TEMP_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011110111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.UN126_TEMP_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_UN123_TEMP_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011110111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.UN123_TEMP_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_UN120_TEMP_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011110111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.UN120_TEMP_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(303),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(302),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(296),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(276),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(272),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(267),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(308),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(271),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(312),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(305),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(299),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(307),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(310),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(309),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_UN132_TEMP_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011110111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.UN132_TEMP_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(280),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(283),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(46),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(269),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(265),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(261),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_COMB_DBGDATA_4_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111001010")
port map (
combout => CPO_DBG_DATAZ(18),
dataa => N_624,
datab => N_688,
datac => N_405,
datad => N_404);
\GRLFPC2_0_COMB_RS2_1_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000010000000")
port map (
combout => \GRLFPC2_0.COMB.RS2_1\(1),
dataa => N_58,
datab => N_17,
datac => \GRLFPC2_0.COMB.RS1_1_SN_M2_I_X\,
datad => \GRLFPC2_0.R.A.RS2\(1));
\GRLFPC2_0_COMB_RS2_1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000010000000")
port map (
combout => \GRLFPC2_0.COMB.RS2_1\(2),
dataa => N_59,
datab => N_17,
datac => \GRLFPC2_0.COMB.RS1_1_SN_M2_I_X\,
datad => \GRLFPC2_0.R.A.RS2\(2));
\GRLFPC2_0_COMB_RS2_1_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000010000000")
port map (
combout => \GRLFPC2_0.COMB.RS2_1\(3),
dataa => N_60,
datab => N_17,
datac => \GRLFPC2_0.COMB.RS1_1_SN_M2_I_X\,
datad => \GRLFPC2_0.R.A.RS2\(3));
\GRLFPC2_0_COMB_RS2_1_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000010000000")
port map (
combout => \GRLFPC2_0.COMB.RS2_1\(4),
dataa => N_61,
datab => N_17,
datac => \GRLFPC2_0.COMB.RS1_1_SN_M2_I_X\,
datad => \GRLFPC2_0.R.A.RS2\(4));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000110000001010")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(12),
dataa => N_618,
datab => N_682,
datac => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datad => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000110000001010")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(15),
dataa => N_621,
datab => N_685,
datac => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datad => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000110000001010")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(19),
dataa => N_625,
datab => N_689,
datac => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datad => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000110000001010")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(20),
dataa => N_626,
datab => N_690,
datac => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datad => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000110000001010")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(21),
dataa => N_627,
datab => N_691,
datac => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datad => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000110000001010")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(28),
dataa => N_634,
datab => N_698,
datac => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datad => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000110000001010")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(29),
dataa => N_635,
datab => N_699,
datac => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datad => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110011111010")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(17),
dataa => N_623,
datab => N_687,
datac => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datad => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110011111010")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(18),
dataa => N_624,
datab => N_688,
datac => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datad => \GRLFPC2_0.COMB.UN1_R.A.RS1_1\);
\GRLFPC2_0_COMB_DBGDATA_4_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111001010")
port map (
combout => CPO_DBG_DATAZ(17),
dataa => N_623,
datab => N_687,
datac => N_405,
datad => N_404);
\GRLFPC2_0_COMB_DBGDATA_4_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011001010")
port map (
combout => CPO_DBG_DATAZ(12),
dataa => N_618,
datab => N_682,
datac => N_405,
datad => N_404);
\GRLFPC2_0_COMB_DBGDATA_4_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011001010")
port map (
combout => CPO_DBG_DATAZ(15),
dataa => N_621,
datab => N_685,
datac => N_405,
datad => N_404);
\GRLFPC2_0_COMB_DBGDATA_4_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011001010")
port map (
combout => CPO_DBG_DATAZ(19),
dataa => N_625,
datab => N_689,
datac => N_405,
datad => N_404);
\GRLFPC2_0_COMB_DBGDATA_4_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011001010")
port map (
combout => CPO_DBG_DATAZ(20),
dataa => N_626,
datab => N_690,
datac => N_405,
datad => N_404);
\GRLFPC2_0_COMB_DBGDATA_4_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011001010")
port map (
combout => CPO_DBG_DATAZ(21),
dataa => N_627,
datab => N_691,
datac => N_405,
datad => N_404);
\GRLFPC2_0_COMB_DBGDATA_4_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011001010")
port map (
combout => CPO_DBG_DATAZ(28),
dataa => N_634,
datab => N_698,
datac => N_405,
datad => N_404);
\GRLFPC2_0_COMB_DBGDATA_4_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011001010")
port map (
combout => CPO_DBG_DATAZ(29),
dataa => N_635,
datab => N_699,
datac => N_405,
datad => N_404);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD55\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(60));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD53\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(61),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(62),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(62),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(63),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(63),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(63),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_64_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(64),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(64),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(64),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_65_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(65),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(65),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_66_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(66),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(66),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(66),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_67_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(67),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(67),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(67),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_68_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(68),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(68),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(68),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_69_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(69),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(69),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(69),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_71_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(71),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(71),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(71),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_72_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(72),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(72),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(72),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_73_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(73),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(73),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(73),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_74_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(74),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(74),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(74),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(75),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(75),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(75),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_76_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(76),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(76),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(76),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_77_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(77),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(77),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_78_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_79_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_80_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(80),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_81_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_82_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(82),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_83_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_84_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD31\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_84_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(84),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD29\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_85_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD30\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_85_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(85),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD28\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_87_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(87),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD28\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(87));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_87_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(87),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD26\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_88_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(88),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD27\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(88));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_88_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(88),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD25\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_89_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(89),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD26\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(89));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_89_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(89),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD24\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_90_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(90),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD25\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(90));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_90_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(90),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD23\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_91_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(91),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD24\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(91));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_91_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(91),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD22\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_92_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(92),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD23\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(92));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_92_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(92),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD21\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_93_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(93),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD22\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(93));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_93_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(93),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD20\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_94_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(94),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD21\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(94));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_94_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(94),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD19\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_95_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(95),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD20\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(95));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_95_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(95),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD18\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_96_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(96),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD19\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(96));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_96_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(96),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD17\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_97_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(97),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD18\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(97));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_97_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(97),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD16\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_99_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(99),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD16\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(99));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_99_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(99),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD14\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_100_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(100),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD15\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(100));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_100_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(100),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD13\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_101_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(101),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD14\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(101));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_101_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(101),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD12\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_102_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(102),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD13\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(102));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_102_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(102),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD11\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_103_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(103),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD12\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(103));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_103_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(103),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD10\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_104_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(104),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD11\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(104));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_104_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(104),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD9\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_105_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(105),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD10\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(105));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_105_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(105),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_106_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(106),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD9\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(106));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_106_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(106),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD7\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_109_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(109),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD6\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(109));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_109_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(109),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_110_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(110),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(110));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_110_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(110),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_111_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(111),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(111));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_111_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(111),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_112_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(112),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(112));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_112_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(112),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_113_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(113),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(113));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_113_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(113),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(26),
dataa => \GRLFPC2_0.R.FSR.TEM\(3),
datab => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datac => \GRLFPC2_0.FPI.OP1_X\(58));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(6),
dataa => \GRLFPC2_0.R.FSR.AEXC\(1),
datab => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datac => \GRLFPC2_0.FPI.OP1_X\(38));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(7),
dataa => \GRLFPC2_0.R.FSR.AEXC\(2),
datab => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datac => \GRLFPC2_0.FPI.OP1_X\(39));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(31),
dataa => \GRLFPC2_0.R.FSR.RD\(1),
datab => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datac => \GRLFPC2_0.FPI.OP1_X\(63));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(30),
dataa => \GRLFPC2_0.R.FSR.RD\(0),
datab => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datac => \GRLFPC2_0.FPI.OP1_X\(62));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(25),
dataa => \GRLFPC2_0.R.FSR.TEM\(2),
datab => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datac => \GRLFPC2_0.FPI.OP1_X\(57));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(24),
dataa => \GRLFPC2_0.R.FSR.TEM\(1),
datab => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datac => \GRLFPC2_0.FPI.OP1_X\(56));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(23),
dataa => \GRLFPC2_0.R.FSR.TEM\(0),
datab => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datac => \GRLFPC2_0.FPI.OP1_X\(55));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(22),
dataa => \GRLFPC2_0.R.FSR.NONSTD\,
datab => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datac => \GRLFPC2_0.FPI.OP1_X\(54));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(14),
dataa => \GRLFPC2_0.R.FSR.FTT\(0),
datab => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datac => \GRLFPC2_0.FPI.OP1_X\(46));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(11),
dataa => CPO_CCZ(1),
datab => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datac => \GRLFPC2_0.FPI.OP1_X\(43));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(10),
dataa => CPO_CCZ(0),
datab => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datac => \GRLFPC2_0.FPI.OP1_X\(42));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(9),
dataa => \GRLFPC2_0.R.FSR.AEXC\(4),
datab => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datac => \GRLFPC2_0.FPI.OP1_X\(41));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(8),
dataa => \GRLFPC2_0.R.FSR.AEXC\(3),
datab => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datac => \GRLFPC2_0.FPI.OP1_X\(40));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(5),
dataa => \GRLFPC2_0.R.FSR.AEXC\(0),
datab => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datac => \GRLFPC2_0.FPI.OP1_X\(37));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(4),
dataa => \GRLFPC2_0.R.FSR.CEXC\(4),
datab => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datac => \GRLFPC2_0.FPI.OP1_X\(36));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(3),
dataa => \GRLFPC2_0.R.FSR.CEXC\(3),
datab => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datac => \GRLFPC2_0.FPI.OP1_X\(35));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(2),
dataa => \GRLFPC2_0.R.FSR.CEXC\(2),
datab => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datac => \GRLFPC2_0.FPI.OP1_X\(34));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(1),
dataa => \GRLFPC2_0.R.FSR.CEXC\(1),
datab => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datac => \GRLFPC2_0.FPI.OP1_X\(33));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(0),
dataa => \GRLFPC2_0.R.FSR.CEXC\(0),
datab => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datac => \GRLFPC2_0.FPI.OP1_X\(32));
\GRLFPC2_0_COMB_RS1_1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.COMB.RS1_1\(2),
dataa => N_84,
datab => \GRLFPC2_0.RS1V_0_SQMUXA_0_A2_X\,
datac => \GRLFPC2_0.COMB.RS1_1_SN_M2_I_X\,
datad => \GRLFPC2_0.COMB.RS1_1_0_X\(2));
\GRLFPC2_0_COMB_RS1_1_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.COMB.RS1_1\(1),
dataa => N_83,
datab => \GRLFPC2_0.RS1V_0_SQMUXA_0_A2_X\,
datac => \GRLFPC2_0.COMB.RS1_1_SN_M2_I_X\,
datad => \GRLFPC2_0.COMB.RS1_1_0_X\(1));
\GRLFPC2_0_COMB_RS1_1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111101101000000")
port map (
combout => \GRLFPC2_0.COMB.RS1_1\(0),
dataa => \GRLFPC2_0.COMB.RS1_1_SN_M2_I_A2\,
datab => N_17,
datac => \GRLFPC2_0.COMB.RS1_1_1_X\(0),
datad => \GRLFPC2_0.COMB.RS1_1_0_X\(0));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(27),
dataa => \GRLFPC2_0.R.FSR.TEM\(4),
datab => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datac => \GRLFPC2_0.FPI.OP1_X\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(20),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(20));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(45),
dataa => N_711,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(161),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(54),
datac => \GRLFPC2_0.FPI.OP2_X\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(51),
datac => \GRLFPC2_0.FPI.OP2_X\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(53),
datac => \GRLFPC2_0.FPI.OP2_X\(50));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(46),
dataa => N_710,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(162),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(52),
datac => \GRLFPC2_0.FPI.OP2_X\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(39),
datac => \GRLFPC2_0.FPI.OP2_X\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(44),
datac => \GRLFPC2_0.FPI.OP2_X\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(21),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(22),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(41),
dataa => N_715,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(157),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(36),
dataa => N_720,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(152),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(24),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(27),
dataa => N_729,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(143),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(35));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(43),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(45),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(45),
datac => \GRLFPC2_0.FPI.OP2_X\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(47),
datac => \GRLFPC2_0.FPI.OP2_X\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(21),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(36),
datac => \GRLFPC2_0.FPI.OP2_X\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(14));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(26),
dataa => N_730,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(142),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(32),
dataa => N_724,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(148),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(41),
datac => \GRLFPC2_0.FPI.OP2_X\(38));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(35),
datac => \GRLFPC2_0.FPI.OP2_X\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(49),
datac => \GRLFPC2_0.FPI.OP2_X\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(50),
dataa => N_706,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(166),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(110));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(53));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(49),
dataa => N_707,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(165),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(52),
dataa => N_704,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(168),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(39),
dataa => N_717,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(155),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(96));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(42),
dataa => N_714,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(158),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(43),
dataa => N_713,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(159),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(37),
dataa => N_719,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(153),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(44),
dataa => N_712,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(160),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(25));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(40),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(40));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(34),
dataa => N_722,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(150),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(33),
dataa => N_723,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(149),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(35),
dataa => N_721,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(151),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(28),
dataa => N_728,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(144),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_41_250_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\(250),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(62),
datac => \GRLFPC2_0.FPI.OP1_X\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_41_252_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\(252),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(60),
datac => \GRLFPC2_0.FPI.OP1_X\(57));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_41_253_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\(253),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(59),
datac => \GRLFPC2_0.FPI.OP1_X\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_41_255_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\(255),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(57),
datac => \GRLFPC2_0.FPI.OP1_X\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_41_256_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\(256),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(53),
datac => \GRLFPC2_0.FPI.OP1_X\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(40),
datac => \GRLFPC2_0.FPI.OP2_X\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_33_244_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_33\(244),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(55),
datac => \GRLFPC2_0.FPI.OP2_X\(52));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_33_238_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_33\(238),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(61),
datac => \GRLFPC2_0.FPI.OP2_X\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(50),
datac => \GRLFPC2_0.FPI.OP2_X\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(51),
datac => \GRLFPC2_0.FPI.OP1_X\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(62),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(53),
datac => \GRLFPC2_0.FPI.OP1_X\(50));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_65_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(65),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(50),
datac => \GRLFPC2_0.FPI.OP1_X\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_68_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(68),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(47),
datac => \GRLFPC2_0.FPI.OP1_X\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_71_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(71),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(44),
datac => \GRLFPC2_0.FPI.OP1_X\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_73_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(73),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(42),
datac => \GRLFPC2_0.FPI.OP1_X\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_74_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(74),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(41),
datac => \GRLFPC2_0.FPI.OP1_X\(38));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_76_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(76),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(39),
datac => \GRLFPC2_0.FPI.OP1_X\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_77_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(77),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(38),
datac => \GRLFPC2_0.FPI.OP1_X\(35));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_79_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(36),
datac => \GRLFPC2_0.FPI.OP1_X\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_80_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(35),
datac => \GRLFPC2_0.FPI.OP1_X\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_245_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\(245),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(232),
datab => NN_2,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD12\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_41_257_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\(257),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(52),
datac => \GRLFPC2_0.FPI.OP1_X\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(46),
datac => \GRLFPC2_0.FPI.OP2_X\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(63),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(52),
datac => \GRLFPC2_0.FPI.OP1_X\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_66_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(66),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(49),
datac => \GRLFPC2_0.FPI.OP1_X\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_69_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(69),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(46),
datac => \GRLFPC2_0.FPI.OP1_X\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(43),
datac => \GRLFPC2_0.FPI.OP2_X\(40));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(37),
datac => \GRLFPC2_0.FPI.OP2_X\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(30),
dataa => N_726,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(146),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111011111000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(38));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(40),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(40));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(40),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(44));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111011111000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(9));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(38));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111011111000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(46),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(41));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(43));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(45),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111011111000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(15));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(16));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(23));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(27));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(31));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(33));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(35));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(36));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(21),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(21));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(21),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(25));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(30));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(14));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(8));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(2),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(1),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(0),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(18));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(20));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(22));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(26));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_A_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10_A\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\(2),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(28),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(28));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(32));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(29),
dataa => N_727,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(145),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(99));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(105));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(112));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(109));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(111));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(88));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(89));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(87));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(91));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(100));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(90));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(92));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(97));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(101));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(102));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(103));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(106));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(21),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(94));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(104));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(93));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(53),
dataa => N_703,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(169),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(40),
dataa => N_716,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(156),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(95));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(31),
dataa => N_725,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(147),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(42),
datac => \GRLFPC2_0.FPI.OP2_X\(39));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_3_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_2\(4));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(46),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(46));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(47),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(47));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(47),
dataa => N_709,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(163),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_41_251_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\(251),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(61),
datac => \GRLFPC2_0.FPI.OP1_X\(58));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_41_254_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_41\(254),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(58),
datac => \GRLFPC2_0.FPI.OP1_X\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_72_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(72),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(43),
datac => \GRLFPC2_0.FPI.OP1_X\(40));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(75),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(40),
datac => \GRLFPC2_0.FPI.OP1_X\(37));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_78_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(37),
datac => \GRLFPC2_0.FPI.OP1_X\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111111100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_33_241_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_33\(241),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(58),
datac => \GRLFPC2_0.FPI.OP2_X\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(50));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_S_8_10_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_S_8_10\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110100001111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_246_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\(246),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD11\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(246));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_251_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\(251),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD6\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(251));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_253_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\(253),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(253));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_255_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\(255),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(255));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_256_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\(256),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(256));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_257_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\(257),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(257));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(372),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_244_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__G1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(244));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_243_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_243__G1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(243));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_242_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_242__G1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(242));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_241_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_241__G1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(241));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_239_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_239__G1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(239));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_237_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_237__G1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(237));
\GRLFPC2_0_COMB_RS1_1_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.COMB.RS1_1\(4),
dataa => N_86,
datab => \GRLFPC2_0.RS1V_0_SQMUXA_0_A2_X\,
datac => \GRLFPC2_0.COMB.RS1_1_SN_M2_I_X\,
datad => \GRLFPC2_0.COMB.RS1_1_0_X\(4));
\GRLFPC2_0_COMB_RS2_1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000010000000")
port map (
combout => \GRLFPC2_0.COMB.RS2_1\(0),
dataa => N_57,
datab => N_17,
datac => \GRLFPC2_0.COMB.RS1_1_SN_M2_I_X\,
datad => \GRLFPC2_0.R.A.RS2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(34));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_64_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(64),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(51),
datac => \GRLFPC2_0.FPI.OP1_X\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111101000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(43),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_3_0_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010111001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_3_0\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(313),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(113),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(17),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(50));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(49));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_108_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(108),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD7\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(108));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_108_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(108),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(108),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_107_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(107),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(107));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_107_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(107),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(107),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD6\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_98_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(98),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD17\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(98));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_98_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(98),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(98),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD15\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP3\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_86_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(86),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD29\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(86));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_A_86_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001111110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_A\(86),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(86),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD27\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP2\,
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNIJE8B_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULTIPLELOGIC_SHIFT_1_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010111001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.MULTIPLELOGIC.SHIFT_1_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(51));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010011000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010011000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010011000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101010100010101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SCTRL_NEW_0_0__G0_I_M2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP2\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD4\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNO_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010111010101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_I_0_0__G0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD5\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(11));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1_REP1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(48),
datac => \GRLFPC2_0.FPI.OP2_X\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(12));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_4_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M2_70_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(70),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(70),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(70),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SS0\);
\GRLFPC2_0_COMB_V_E_STDATA_1_1_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(16),
dataa => \GRLFPC2_0.R.FSR.FTT\(2),
datab => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datac => \GRLFPC2_0.FPI.OP1_X\(48));
\GRLFPC2_0_COMB_V_E_STDATA_1_1_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111100100000")
port map (
combout => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(13),
dataa => \GRLFPC2_0.R.STATE\(1),
datab => \GRLFPC2_0.R.STATE\(0),
datac => \GRLFPC2_0.COMB.V.A.AFSR_1\,
datad => \GRLFPC2_0.FPI.OP1_X\(45));
\GRLFPC2_0_COMB_DBGDATA_4_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010011100100")
port map (
combout => CPO_DBG_DATAZ(13),
dataa => N_404,
datab => \GRLFPC2_0.COMB.DBGDATA_4_0_X\(13),
datac => \GRLFPC2_0.R.STATE\(1),
datad => \GRLFPC2_0.R.STATE\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_67_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(67),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(48),
datac => \GRLFPC2_0.FPI.OP1_X\(45));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_19_70_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(70),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP1_X\(45),
datac => \GRLFPC2_0.FPI.OP1_X\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(38),
dataa => N_718,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(154),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_250_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\(250),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD7\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(250));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_248_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\(248),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD9\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(248));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_247_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\(247),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD10\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(247));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_33_242_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_33\(242),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(57),
datac => \GRLFPC2_0.FPI.OP2_X\(54));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_249_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\(249),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(249));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_33_239_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_33\(239),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(60),
datac => \GRLFPC2_0.FPI.OP2_X\(57));
GRLFPC2_0_COMB_FPDECODE_RS1D5_0_A2_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000010000")
port map (
combout => \GRLFPC2_0.COMB.FPDECODE.RS1D5_0_A2_0\,
dataa => N_69,
datab => N_70,
datac => N_63,
datad => N_62);
\GRLFPC2_0_COMB_RS1_1_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC2_0.COMB.RS1_1\(3),
dataa => N_85,
datab => \GRLFPC2_0.RS1V_0_SQMUXA_0_A2_X\,
datac => \GRLFPC2_0.COMB.RS1_1_SN_M2_I_X\,
datad => \GRLFPC2_0.COMB.RS1_1_0_X\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_33_240_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_33\(240),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(59),
datac => \GRLFPC2_0.FPI.OP2_X\(56));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_33_237_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_33\(237),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(62),
datac => \GRLFPC2_0.FPI.OP2_X\(59));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_238_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_238__G1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(238));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNO_0_240_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_240__G1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(240));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_254_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\(254),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(254));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2_252_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_2\(252),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(252));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_33_243_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_33\(243),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(56),
datac => \GRLFPC2_0.FPI.OP2_X\(53));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_11_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011110000111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_11_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(48),
dataa => N_708,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(164),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(51),
dataa => N_705,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(167),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_1_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_1\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.OP2_X\(38),
datac => \GRLFPC2_0.FPI.OP2_X\(35));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_3_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_3\(54),
dataa => N_702,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(170),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datad => \GRLFPC2_0.FPI.LDOP_REP3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(277),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(0),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_14_2_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_14_2\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_1162\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_12_0_A2\(62));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110000001100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_12\(60));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_12\(60));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_11_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_11\(62),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_1_0_A2_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_1_0_A2\(62),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_2_0_A2_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_2_0_A2\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_36_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_36\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_A26_17_0_A2_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_A26_17_0_A2\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_10_1_0_A2_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_10_1_0_A2\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_37_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_37\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_8_RNIJMU96: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_4785_A2_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_8_RNIJMU96_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_4859_A2_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_11_0_A2_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_11_0_A2\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_35_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_35\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_RNO_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_4510_A2_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_0_A2_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_0_A2\(46),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_25_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_25\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111101111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_0_I_O2_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_O2\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_0_I_O2_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_0_I_O2\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A26_2_0_I_O2_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A26_2_0_I_O2\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_12_I_O2_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111101111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_12_I_O2\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_6_I_O2_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111111011111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_6_I_O2\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_17_1_I_O2_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111110111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_17_1_I_O2\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A2_3_I_O2_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111110111111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_3_I_O2\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O20_3_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100011111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O20_3\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_19_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_19\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O16_0_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101111001011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_0\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_X2_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101100101011001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O23_5_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101010111010101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_5\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A2_7_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010011000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A2_7\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_O28_1_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010001110100011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_O28_1\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_O2_3_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011110010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_O2_3\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O26_5_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100011111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O26_5\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_9_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000001010000010")
port map (
combout => NN_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O22_9_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110111001101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_9\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_4_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_4\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_5_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_5\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A2_9_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A2_9\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_M27_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111110001111100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_M27\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_X2_0_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101011001010110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_X2_0\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_O27_2_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111011111110111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_O27_2\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_7_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010000010100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_7\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_8_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O22_3_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000110110001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_3\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O22_5_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101011000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_5\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_X2_2_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101011001010110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_X2_2\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_1_M24_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111010011110000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_1_M24\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_O23_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110110001101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O23\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_5_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_5\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_11_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_11\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O27_10_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O27_10\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_6_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100110001001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_6\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_1_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_1\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_O30_7_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101110101111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_O30_7\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_3_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110010001100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O21_2_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O21_2\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O21_3_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101110101011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O21_3\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_5_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_5\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_M2_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101000111100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_M2\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O28_5_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110011101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O28_5\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_M2_0_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011010000110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_M2_0\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_I_O2_2_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000101110001011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_O2_2\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_8_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_18_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_18\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_20_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_20\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_M2_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011010000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_M2\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_5_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_5\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O18_6_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O18_6\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O20_6_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O20_6\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_8_RNIVFEF3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_9_7495\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_5_1_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000101000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_5_1\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_7_2_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7_2\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_11_2_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11_2\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_13_2_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001000010010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_13_2\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_14_2_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001000010010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_14_2\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_17_1_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_17_1\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_18_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_18\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_1_0\(5));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_10_1_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_10_1\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_25_1_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_25_1\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A29_22_1_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A29_22_1\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_7_1_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010100010101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_7_1\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_11_1_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101010001010100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11_1\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_12_2_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_12_2\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_17_1_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_17_1\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_20_4_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_20_4\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_26_2_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_26_2\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_34_2_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_34_2\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_1_2_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_1_2\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_2_3_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_2_3\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A15_11_2_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_11_2\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_8_2_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_8_2\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_16_1_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_16_1\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_18_3_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_18_3\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_A27_20_2_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_A27_20_2\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_2_2_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_2_2\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_13_2_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_13_2\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_16_2_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_16_2\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_5_1_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_5_1\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_6_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_6\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A24_10_1_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_10_1\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A24_17_2_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_17_2\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A24_18_1_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_18_1\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A24_20_2_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_20_2\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_8_1_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_8_1\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_14_3_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_14_3\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_13_1_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_13_1\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_24_3_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_24_3\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A19_2_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A19_2\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_0_2_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_0_2\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_4_2_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_4_2\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_13_1_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_13_1\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_21_2_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_21_2\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A30_12_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_12\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A30_15_2_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_15_2\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_I_A30_26_2_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_I_A30_26_2\(60),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A21_1_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001000010010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A21_1\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_1_1_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_1_1\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_2_2_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_2_2\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_16_2_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_16_2\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_18_2_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_18_2\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_2_2_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_2_2\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_18_3_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_18_3\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_22_1_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_22_1\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_I_I_A26_1_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_I_A26_1\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_1_0_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_1_0\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_0_2_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_0_2\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A21_2_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A21_2\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_4_4_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_4\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_15_3_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_15_3\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_15_4_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_15_4\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_7_2_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_7_2\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_12_2_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_12_2\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_13_1_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_13_1\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A7_2_4_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A7_2_4\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A3_3_2_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A3_3_2\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_0_2_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_2\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_5_4_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_4\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_2_1_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_2_1\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_1_2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001000010010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_1_2\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_2_1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_2_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_4_2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_4_2\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_5_3_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_5_3\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_1_2_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_1_2\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_0_1_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => N_34483_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_I_A26_6_1_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_I_I_A26_6_1\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_7_2_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_7_2\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_4_1_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_1\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_11_4_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_4\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_6_2_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_6_2\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_5_1_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_5_1\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_A24_0_2_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_A24_0_2\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(83),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_2_0_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_2_0\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_1_A2_1_1_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1_A2_1_1\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_1_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0_1\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_4_1_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_4_1\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101000001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_1\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_16_4_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_16_4\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datad => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_25_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_4_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_C\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGXZ_UN5_XZAREGLOADEN_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLAREGXZ.UN5_XZAREGLOADEN_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNI754D_77_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW_0\(77),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN13_INEXACT_9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.INEXACTSIG.UN13_INEXACT_9\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30));
GRLFPC2_0_COMB_V_A_AFQ_1_4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.COMB.V.A.AFQ_1_4\,
dataa => \GRLFPC2_0.R.A.ST_RET_2\(1),
datab => \GRLFPC2_0.R.A.AFQ_RET\(9));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN7_FEEDBACK_0_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN7_FEEDBACK_0_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(51));
GRLFPC2_0_COMB_UN2_HOLDN_0_A2_11_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_11_0\,
dataa => \GRLFPC2_0.R.A.MOV_RET\(9),
datab => \GRLFPC2_0.R.A.MOV_RET\(13));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_RESULT_U_RNO_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111011101110111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.G_31_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(50));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN1_S_DYADIC_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN1_S_DYADIC_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN7_FEEDBACK_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.FEEDBACKMULXFF.UN7_FEEDBACK_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(49));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN6_U_RDN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.UN6_U_RDN\,
dataa => \GRLFPC2_0.R.FSR.RD\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(198),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(189),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(188),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(176),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP3\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPYBUS_2_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(316),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(341),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(338),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(337),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(214),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(46),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(185),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(178),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(195),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(40),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(191),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(40),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(184),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(46),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(205),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(190),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(174),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110111011101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110111011101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110111011101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(21),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(210),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(206),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(199),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(192),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(175),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(177),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_XZBREGLC_2_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLBREGXZ.XZBREGLC_2\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
datab => \GRLFPC2_0.FPI.LDOP_REP0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGXZ_UN4_XZBREGLOADEN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLBREGXZ.UN4_XZBREGLOADEN\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_V_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELECTQUOBITS_NOTDIVC_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.SELECTQUOBITS.NOTDIVC\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(375),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(374));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RNISH49_376_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.SELECTQUOBITS.NOTDIVC\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(376),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(374));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(212),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(211),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(17));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(347),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(346),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(345),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(344),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(343),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(342),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(340),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(339),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(336),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(335),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(334),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(40),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(333),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(368),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(367),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(366),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(365),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(364),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(363),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(362),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(361),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(360),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(359),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(358),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(357),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(356),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(355),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(354),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(353),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(21),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(352),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(351),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(350),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(349),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(348),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(324),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(326),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(325),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(323),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(322),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(321),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(320),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(319),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(318),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(317),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(332),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(331),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(330),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(329),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(45),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(328),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(46),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(327),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(200),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(213),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(209),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(208),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(207),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(204),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(203),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(202),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(193),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(196),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_ROMXZSL2FROMC: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.ROMXZSL2FROMC\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(194),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD56\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(61),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD54\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(62),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD53\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(63),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(63),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD52\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_64_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(64),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(64),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD51\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_65_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(65),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD50\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_66_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(66),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD49\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_67_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(67),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(67),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD48\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_68_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(68),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(68),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD47\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_69_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(69),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(69),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD46\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_71_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(71),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(71),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD44\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_72_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(72),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(72),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD43\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_73_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(73),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(73),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD42\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_74_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(74),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(74),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD41\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(75),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(75),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD40\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_76_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(76),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(76),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD39\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_77_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(77),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD38\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_78_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD37\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_79_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD36\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_80_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD35\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_81_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD34\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_82_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD33\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_83_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD32\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_114_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(114),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD52\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(62),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD51\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(63),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD50\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_64_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(64),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD49\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_65_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(65),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD48\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_66_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(66),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD47\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_67_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(67),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD46\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_68_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(68),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD45\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_69_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(69),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD44\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_71_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(71),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD42\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_72_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(72),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD41\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_73_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(73),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD40\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_74_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(74),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD39\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(75),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD38\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_76_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(76),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD37\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_77_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(77),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD36\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_78_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(78),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD35\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_79_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(79),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD34\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_80_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(80),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD33\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_81_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(81),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD32\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_82_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(82),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD31\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_83_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(83),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD30\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\);
\GRLFPC2_0_COMB_V_I_PC_1_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(22),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(20),
datab => \GRLFPC2_0.R.I.PC_RET\(20),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(8),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(6),
datab => \GRLFPC2_0.R.I.PC_RET\(6),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(7),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(5),
datab => \GRLFPC2_0.R.I.PC_RET\(5),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(12),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(10),
datab => \GRLFPC2_0.R.I.PC_RET\(10),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(11),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(9),
datab => \GRLFPC2_0.R.I.PC_RET\(9),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(10),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(8),
datab => \GRLFPC2_0.R.I.PC_RET\(8),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(9),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(7),
datab => \GRLFPC2_0.R.I.PC_RET\(7),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(16),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(14),
datab => \GRLFPC2_0.R.I.PC_RET\(14),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(15),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(13),
datab => \GRLFPC2_0.R.I.PC_RET\(13),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(14),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(12),
datab => \GRLFPC2_0.R.I.PC_RET\(12),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(13),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(11),
datab => \GRLFPC2_0.R.I.PC_RET\(11),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(21),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(19),
datab => \GRLFPC2_0.R.I.PC_RET\(19),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(20),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(18),
datab => \GRLFPC2_0.R.I.PC_RET\(18),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(31),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(29),
datab => \GRLFPC2_0.R.I.PC_RET\(29),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(30),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(28),
datab => \GRLFPC2_0.R.I.PC_RET\(28),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(27),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(25),
datab => \GRLFPC2_0.R.I.PC_RET\(25),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(26),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(24),
datab => \GRLFPC2_0.R.I.PC_RET\(24),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(29),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(27),
datab => \GRLFPC2_0.R.I.PC_RET\(27),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(25),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(23),
datab => \GRLFPC2_0.R.I.PC_RET\(23),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(18),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(16),
datab => \GRLFPC2_0.R.I.PC_RET\(16),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(17),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(15),
datab => \GRLFPC2_0.R.I.PC_RET\(15),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(28),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(26),
datab => \GRLFPC2_0.R.I.PC_RET\(26),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(6),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(4),
datab => \GRLFPC2_0.R.I.PC_RET\(4),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(5),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(3),
datab => \GRLFPC2_0.R.I.PC_RET\(3),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(4),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(2),
datab => \GRLFPC2_0.R.I.PC_RET\(2),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(3),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(1),
datab => \GRLFPC2_0.R.I.PC_RET\(1),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(2),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(0),
datab => \GRLFPC2_0.R.I.PC_RET\(0),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(24),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(22),
datab => \GRLFPC2_0.R.I.PC_RET\(22),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_COMB_V_I_PC_1_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(23),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(21),
datab => \GRLFPC2_0.R.I.PC_RET\(21),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD37\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD38\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(20),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD36\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD37\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD33\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD34\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD29\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD30\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD48\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD49\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD47\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD48\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD54\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD55\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD49\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD50\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD52\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD53\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(21),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(21),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD35\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD36\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(22),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD34\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD35\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD2\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD17\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD18\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD32\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD33\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(45),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD25\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD26\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD21\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD22\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD15\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD16\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD13\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD14\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(45),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD11\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD12\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(26),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD30\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD31\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD43\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD44\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD41\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD42\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(16),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD40\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD41\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(14),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD42\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD43\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000110110001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD57\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD20\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD21\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD1\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD4\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD5\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD12\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD13\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD8\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD9\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD3\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD4\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD14\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD15\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(37),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD19\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD20\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(21),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD31\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD32\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(40),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(40),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD16\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD17\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_118_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_118\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(18),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(17),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(60));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD39\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD40\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD38\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD39\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_235_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(235),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD9\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_239_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(239),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(252),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD5\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_243_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(243),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(256),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_244_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(244),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(257),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD51\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD52\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_MIXOIN_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.MIXOIN\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(35),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_2\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(257),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_237_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(237),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(250),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD7\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD23\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD24\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_233_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(233),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD11\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD18\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD19\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100110101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(46),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD27\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD28\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD26\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD27\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(17),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(238),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(239),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(240),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(2),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(41),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(241),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(35),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(23),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(15),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(28),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD28\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD29\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(32),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD24\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD25\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD56\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD57\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_2\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(251),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(238));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_2\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(252),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(239));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_2\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(253),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(240));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_0_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.EXPYBUS_0\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(240));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD53\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD54\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_2\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(250),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(237));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(46),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(46),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD10\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD11\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD9\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD10\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_241_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(241),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(254),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_246_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(246),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD12\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_251_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(251),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(238),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD7\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_253_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(253),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(240),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD5\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_255_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(255),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_256_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(256),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_257_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(257),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_242_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(242),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(255),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TOPBITSIN\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(237),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_SUB_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110110001101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(19));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(1),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD55\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD56\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DECODESTATUS_UN7_STATUS: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DECODESTATUS.UN7_STATUS\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(39),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(38));
GRLFPC2_0_COMB_V_A_AFSR_1_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.COMB.V.A.AFSR_1_2\,
dataa => \GRLFPC2_0.R.A.MOV_RET\(15),
datab => \GRLFPC2_0.R.A.AFQ_RET\(5));
GRLFPC2_0_COMB_V_A_AFSR_1_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.N_782\,
dataa => \GRLFPC2_0.R.A.AFQ_RET\(9),
datab => \GRLFPC2_0.R.A.MOV_RET\(0));
GRLFPC2_0_COMB_QNE2_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.COMB.QNE2_0\,
dataa => \GRLFPC2_0.R.A.SEQERR_RET_4\(0),
datab => \GRLFPC2_0.R.A.SEQERR_RET_4\(1));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPAREGLOADEN_RNICN17: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101110111011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M2_0\,
dataa => \GRLFPC2_0.FPI.LDOP_REP5\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPAREGLOADEN\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD22\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD23\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_ADD3\);
GRLFPC2_0_FPCO_HOLDN_0_I: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => CPO_HOLDNZ,
dataa => \GRLFPC2_0.R.MK.BUSY_RET_5\,
datab => \GRLFPC2_0.R.MK.HOLDN2\);
GRLFPC2_0_COMB_UN6_IUEXEC_RNIBU97: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => G_8482,
dataa => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2\,
datab => \GRLFPC2_0.COMB.UN6_IUEXEC\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_REP4_RNI65S9_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIDVK7_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111011101110111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_AREGXORBREG_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SFTLFT.AREGXORBREG_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN1_GRFPUS: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SFTLFT.UN1_GRFPUS\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(24));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(179),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(197),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(42),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_116_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_116\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(10),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD50\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD51\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(181),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(182),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD6\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD7\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(50),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD7\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD8\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIGOP2_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(5),
datab => \GRLFPC2_0.FPI.LDOP_REP5\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(373),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(0));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_0_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_0\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(10));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD5\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD6\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(46),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.TEMP\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD45\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD46\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(11),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(43),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD44\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD45\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(12),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.RIGHTSHIFTERBL.S_8\(45),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SRCONTROL_1\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_1_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_1\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD46\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD47\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_2_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_2\(10),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_ADD3\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M1_70_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M1\(70),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD43\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_70_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(70),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD45\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(45),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(70));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(45),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(186),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2_REP1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_TEMP_1_1_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(187),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2_REP1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN1_TEMP: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN1_TEMP\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(72));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNO_74_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_74__G0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(62),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT\);
\GRLFPC2_0_COMB_V_I_PC_1_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC2_0.COMB.V.I.PC_1\(19),
dataa => \GRLFPC2_0.R.I.PC_RET_30\(17),
datab => \GRLFPC2_0.R.I.PC_RET\(17),
datac => \GRLFPC2_0.R.I.PC_RET_60\);
GRLFPC2_0_COMB_PEXC8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => CPO_EXCZ,
dataa => \GRLFPC2_0.R.STATE\(1),
datab => \GRLFPC2_0.R.STATE\(0));
\GRLFPC2_0_R_STATE_RNI9D7D_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.N_1213_I_0_O2\,
dataa => \GRLFPC2_0.R.STATE\(0),
datab => \GRLFPC2_0.R.STATE\(1));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.S_8\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_250_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(250),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(237),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD8\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_248_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(248),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD10\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_247_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(247),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD11\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_2\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(249),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS_2_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_2\(9),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_249_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(249),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD9\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_236_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(236),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(249),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD8\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => NN_2,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RNIQ83D_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_SN_M3_E\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(43),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_EXPBREGLOADEN_RNIDN17: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101110111011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_1\,
dataa => \GRLFPC2_0.FPI.LDOP_REP5\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_234_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(234),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(247),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD10\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_254_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(254),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(241),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD4\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_252_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(252),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(239),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD6\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_238_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(238),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(251),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD6\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_232_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(232),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(245),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD12\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_240_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1\(240),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(253),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD4\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_17: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_17\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD56\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD57\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_M0_115_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M0\(115),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(115),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD0\,
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2S2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_9_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001100110011001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_9_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_8_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001100110011001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_8_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RNIRH78_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111011101110111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
datab => \GRLFPC2_0.FPI.LDOP_REP0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(38),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(77));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_1_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_1\(24),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_11_2\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A2_9_0_A2\(61));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_1_A2_3_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_1_A2_3\(39),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_4785_A2_2\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_O12_0_A2_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_O12_0_A2\(44),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_18_2\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A15_3_1\(18));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_8_RNI2AOD3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8577_I_0_A2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_12_RNI42TE3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_8466_I_I_I_X2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_1_0_A2_RNO_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_11846_I_I_I_X2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_X2_0_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_0\(30),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A2_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_X2_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(29),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_X2_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_M2_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101000111010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_M2\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_M2_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_M2\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_M29_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000101110001011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_M29\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A2_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_X2_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_M23_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000101110001011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_M23\(52),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_0_O28_5_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101110111011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_O28_5\(56),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A2_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_X2_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_X2\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_M26_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_M26\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_X2_0_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_0\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_M22_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_M22\(53),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A2_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_I_I_I_0_M27_0_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0_M27_0\(47),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_X2_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_O25_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110111011101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O25\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_X2_1_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_1\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_M2_0_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000101110001011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_M2_0\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O22_1_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111011101110111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O22_1\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_M2_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000110110001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_M2\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_M2_0_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101000111010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_M2_0\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_X2_0_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_0\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_8_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_X2_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_O2_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101110111011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O2\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O23_1_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111011101110111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O23_1\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_M2_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_M2\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_3_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A2_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A2\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O19_1_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111011101110111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_1\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O19_2_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110111011101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_8_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_3_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_3\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_5_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_5\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_M21_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_M21\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_2_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_2\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_X2_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O2_2_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111011101110111")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O2_2\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_I_I_X2_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_I_I_X2\(31),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_O21_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101110111011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O21\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_X2_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_X2_3_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_3\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_X2_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_X2_0_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_0\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_M17_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_M17\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A3_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A3\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_X3_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X3\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O16_0_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110111011101")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O16_0\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_X2_0_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_X2_0\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_M16_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_M16\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78),
datac => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_0_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_0\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A2_8_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A2_8\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_O18_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O18\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O18_4_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O18_4\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A2\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O13_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O13_0\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_X2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_X2\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_A12_0_I_2_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101110111011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_A12_0_I_2\(25),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A14_1_1_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A14_1_1\(62),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_0_1_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_1\(49),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A23_1_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(33),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A29_1_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\(58),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A26_1_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A26_1\(55),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A15_1_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A15_1\(18),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A25_1_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A25_1\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_16_1_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A25_16_1\(27),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A22_1_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A22_1\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_4_2_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_4_2\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_12_1_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_12_1\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_13_1_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_13_1\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_17_1_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => N_33157_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_9_1_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_9_1\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A23_14_2_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A23_14_2\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A27_16_1_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A27_16_1\(54),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A19_1_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A19_1\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_4_1_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_4_1\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_6_1_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_6_1\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A19_14_1_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A19_14_1\(13),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A13_1_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A13_1\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_0_1_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_0_1\(48),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A28_1_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A28_1\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A28_12_1_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A28_12_1\(57),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_I_I_A26_20_1_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => N_34381_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_2_1_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_2_1\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_3_1_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_3_1\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A20_5_1_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A20_5_1\(36),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_4_1_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_1\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_4_2_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_4_2\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_7_1_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => N_33227_2,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_16_1_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_16_1\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A17_1_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A17_1\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_3_1_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => N_28709_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_7_1_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_7_1\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A17_8_1_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A17_8_1\(34),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A7_1_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A7_1\(3),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_1_0_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => N_34072_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_0_1_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_0_1\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_2_1_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_2_1\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_3_1_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_3_1\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_4_1_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_4_1\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_5_1_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_1\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_5_2_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_5_2\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_11_1_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => N_29496_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_11_2_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_11_2\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_12_1_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_12_1\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A16_13_1_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A16_13_1\(5),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_3_1_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => N_28871_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_7_1_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_7_1\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_8_1_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_8_1\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_9_1_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_9_1\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_10_1_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_10_1\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_13_1_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_13_1\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A18_14_1_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A18_14_1\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A13_1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A13_2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A13_2\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_1_1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_1_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_5_1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_5_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_7_1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_7_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(84));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_9_1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_9_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_10_1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_10_1\(0),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(81));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A21_1_1_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A21_1_1\(51),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_11_1_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_1\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_11_2_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_11_2\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(78),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_5_1_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_5_1\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(80));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A22_1_1_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A22_1_1\(6),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_1_A29_1_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_1_A29_1\(19),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN3_S_SQRT_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => N_33495_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(78));
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN3_S_SQRT_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.ENTRYSHFT.UN3_S_SQRT_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A13_16_2_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_16_2\(61),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(78));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_A23_1_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_A23_1\(59),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(81),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_A25_7_1_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => N_32980_1,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(79));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_0_O2_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101110111011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_0_O2\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(83));
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_0_O18_0_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101110111011")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O18_0\(4),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP5\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP6\(80));
GRLFPC2_0_R_M_AFSR_RET_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.R.M.AFSR_RET_0_0_G1\,
dataa => \GRLFPC2_0.R.E.AFSR_RET\,
datab => \GRLFPC2_0.R.E.AFQ_RET_1\);
GRLFPC2_0_R_M_AFQ_RET_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC2_0.R.M.AFQ_RET_0_0_G1\,
dataa => \GRLFPC2_0.R.E.AFQ_RET\,
datab => \GRLFPC2_0.R.E.AFQ_RET_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_ADD12: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011010010110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD12\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(12),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(12),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_11\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_ADD11: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD11\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_11\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(11),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_10\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_ADD10: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD10\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_10\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(10),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_9\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_ADD9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD9\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_9\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(9),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_8\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_ADD8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD8\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_8\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(8),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_7\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_ADD7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD7\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(7),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_6\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_ADD6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD6\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_6\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(6),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_5\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_ADD5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD5\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_5\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(5),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_4\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_ADD4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD4\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(4),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_ADD3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD3\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_ADD2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_ADD1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_ADD0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPXBUS_3\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_V_0\(0),
cin => N_58394);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD57: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011010010110")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD57\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(57),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(57),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_56\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD56: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD56\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_56\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(56),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(56),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_55\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD55: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD55\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_55\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(55),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(55),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_54\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD54: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD54\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_54\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(54),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(54),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_53\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD53: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD53\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_53\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(53),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(53),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_52\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD52: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD52\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_52\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(52),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(52),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_51\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD51: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD51\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_51\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(51),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(51),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_50\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD50: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD50\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_50\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(50),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(50),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_49\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD49: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD49\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_49\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(49),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(49),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_48\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD48: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD48\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_48\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(48),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(48),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_47\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD47: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD47\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_47\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(47),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(47),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_46\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD46: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD46\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_46\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(46),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(46),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_45\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD45: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD45\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_45\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(45),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(45),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_44\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD44: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD44\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_44\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(44),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(44),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_43\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD43: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD43\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_43\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(43),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(43),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_42\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD42: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD42\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_42\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(42),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(42),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_41\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD41: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD41\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_41\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(41),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(41),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_40\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD40: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD40\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_40\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(40),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(40),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_39\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD39: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD39\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_39\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(39),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(39),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_38\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD38: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD38\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_38\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(38),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(38),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_37\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD37: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD37\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_37\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(37),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(37),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_36\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD36: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD36\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_36\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(36),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(36),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_35\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD35: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD35\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_35\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(35),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(35),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_34\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD34: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD34\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_34\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(34),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(34),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_33\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD33: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD33\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_33\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(33),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(33),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_32\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD32: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD32\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_32\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(32),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(32),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_31\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD31: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD31\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_31\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(31),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(31),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_30\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD30: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD30\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_30\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(30),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(30),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_29\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD29: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD29\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_29\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(29),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(29),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_28\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD28: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD28\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_28\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(28),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(28),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_27\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD27: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD27\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_27\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(27),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(27),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_26\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD26: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD26\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_26\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(26),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(26),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_25\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD25: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD25\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_25\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(25),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(25),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_24\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD24: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD24\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_24\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(24),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(24),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_23\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD23: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD23\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_23\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(23),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(23),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_22\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD22: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD22\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_22\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(22),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(22),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_21\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD21: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD21\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_21\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(21),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(21),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_20\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD20: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD20\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_20\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(20),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(20),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_19\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD19: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD19\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_19\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(19),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(19),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_18\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD18: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD18\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_18\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(18),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(18),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_17\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD17: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD17\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_17\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(17),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(17),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_16\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD16: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD16\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_16\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(16),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(16),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_15\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD15: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD15\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_15\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(15),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(15),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_14\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD14: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD14\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_14\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(14),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(14),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_13\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD13: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD13\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_13\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(13),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(13),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_12\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD12: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD12\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_12\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(12),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(12),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_11\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD11: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD11\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_11\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(11),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(11),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_10\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD10: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD10\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_10\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(10),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(10),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_9\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD9\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_9\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(9),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(9),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_8\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD8\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_8\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(8),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(8),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_7\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD7\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(7),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(7),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_6\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD6\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_6\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(6),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(6),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_5\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD5\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_5\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(5),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(5),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_4\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD4\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(4),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(4),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100110110010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD3\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(3),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_3_M4_I_X2\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(2),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(1),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF_ADD0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0\(0),
cin => N_58395);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_PCTRL_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0101101001011010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL\(8),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(78),
datab => GND,
cin => N_30136);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_PCTRL_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110110001101100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL\(7),
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
cin => N_30135);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_PCTRL_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0101101010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL\(6),
cout => N_30136,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(80),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(79),
cin => N_30134);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_PCTRL_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110110010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL\(5),
cout => N_30135,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
cin => N_30133);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_PCTRL_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0101101010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL\(4),
cout => N_30134,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP7\(82),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(81),
cin => N_30132);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_PCTRL_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110110010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL\(3),
cout => N_30133,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83),
cin => N_30130);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_PCTRL_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0101101010000000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL\(2),
cout => N_30132,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(84),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(83),
cin => N_30129);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_PCTRL_A_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000000100010")
port map (
cout => N_30129,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_PCTRL_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001100100100010")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL\(1),
cout => N_30130,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP8\(85),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_ADD12: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100101101001")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD12\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(232),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(245),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_11\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_ADD11: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD11\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_11\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_10\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_ADD10: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD10\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_10\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(247),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_9\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_ADD9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD9\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_9\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_8\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_ADD8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD8\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_8\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(249),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_7\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_ADD7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD7\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_7\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(237),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(250),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_6\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_ADD6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD6\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_6\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(238),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(251),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_5\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_ADD5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD5\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_5\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(239),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(252),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_4\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_ADD4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD4\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_4\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(240),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(253),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_3\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_ADD3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD3\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_3\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(241),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(254),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_ADD2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(255),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_ADD1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(256),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_0\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_ADD0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.GRFPUE_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(257),
cin => N_58396);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_3_RNID2884: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_ADD3\,
cout => N_58397,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_2_RNIEF0T1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIHA5S_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI7NQB_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(34),
cin => N_58398);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_1_RNI7NR24: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_ADD3\,
cout => N_58399,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_RNICJ712: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_1_RNIPRNR: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI8NQ8_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(33),
cin => N_58400);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_3_RNIVFBG3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_ADD3\,
cout => N_58401,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_60_SUM1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_RNIS16M1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_60_SUM0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIFT0U_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.CI_2_SUM0_0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI5FBE_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57),
cin => N_58402);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_3_RNI345R3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_ADD3\,
cout => N_58403,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_1_RNID8212: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_RNISQRR: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI8BVA_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(56),
cin => N_58404);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_2_RNI7CTR3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_ADD3\,
cout => N_58405,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_RNIFBIO1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIMDMP_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIA7J7_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(55),
cin => N_58406);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_RNI7CCO3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_ADD3\,
cout => N_58407,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_RNI3ACM1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI06IN_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIE37C_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(54),
cin => N_58408);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_3_RNIGKEF3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_ADD3\,
cout => N_58409,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_3_RNINHHL1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_1_RNINS5N: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIGVQ8_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(53),
cin => N_58410);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_3_RNIT93F3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_ADD3\,
cout => N_58411,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_2_RNIBVCH1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIGJPM_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI2Q67_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(52),
cin => N_58412);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_RNI77NC3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_ADD3\,
cout => N_58413,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_2_RNI2D8L1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI9ADM_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI4MQB_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(51),
cin => N_58414);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_3_RNI9N4O3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_ADD3\,
cout => N_58415,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_3_RNI2HFP1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIANCU_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIU6IA_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(50),
cin => N_58416);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_1_RNIMG654: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_ADD3\,
cout => N_58417,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_2_RNIC6M52: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIFVVT_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI3UPE_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(49),
cin => N_58418);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_1_RNI0FT64: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_ADD3\,
cout => N_58419,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_3_RNI7FIU1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_RNIVVKQ: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNISEN9_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(48),
cin => N_58420);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_RNI4CDF4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_ADD3\,
cout => N_58421,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_3_RNIALM72: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI37KV_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIVRMC_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(19),
cin => N_58422);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_1_RNI2KVP4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_ADD3\,
cout => N_58423,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_2_RNIJ9HE2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_RNIGSKA1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI1QRM_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(18),
cin => N_58424);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_3_RNIBD014: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_ADD3\,
cout => N_58425,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_3_RNIG45R1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIJKUT_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIVABE_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(47),
cin => N_58426);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_3_RNIC4G04: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_ADD3\,
cout => N_58427,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_1_RNI36E12: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_RNIF1AS: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI2MDB_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(46),
cin => N_58428);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_2_RNIF0JT3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_ADD3\,
cout => N_58429,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_1_RNI22SP1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIDGOP_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI63J7_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(45),
cin => N_58430);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_2_RNICN8K3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_ADD3\,
cout => N_58431,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_1_RNIRSFJ1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIMTHN_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI9V6C_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(44),
cin => N_58432);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_RNIVTRD3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_ADD3\,
cout => N_58433,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_3_RNIPJNK1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_3_RNI47CM: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI1E18_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(43),
cin => N_58434);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_2_RNIB65I3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_ADD3\,
cout => N_58435,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_1_RNIPP8L1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIJ3FR_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIFT4A_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(42),
cin => N_58436);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_RNIUG6O3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_ADD3\,
cout => N_58437,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_3_RNICSRS1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIG9BP_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIUHQB_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(41),
cin => N_58438);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_1_RNII8I04: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_ADD3\,
cout => N_58439,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_1_RNI4J9Q1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI8Q8S_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI3EE8_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(40),
cin => N_58440);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_RNI003R3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_ADD3\,
cout => N_58441,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_RNIL4AQ1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIE2SR_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIUPPE_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(39),
cin => N_58442);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_1_RNI9BK14: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_ADD3\,
cout => N_58443,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_1_RNIDHI32: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI9VO11_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIPAN9_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(38),
cin => N_58444);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_2_RNIC27E4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_ADD3\,
cout => N_58445,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_2_RNIIR822: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIDCUT_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIS6BE_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(37),
cin => N_58446);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_RNIGOBC4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_ADD3\,
cout => N_58447,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_1_RNINKS52: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_3_RNIAOO01: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIU2VA_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(36),
cin => N_58448);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_3_RNIH7GC4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_ADD3\,
cout => N_58449,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_2_RNILU732: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI5MLU_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNII4K7_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(35),
cin => N_58450);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_1_RNIPUJ24: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_ADD3\,
cout => N_58451,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_2_RNIUS7V1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIP9KU_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI3E1B_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(7),
cin => N_58452);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_2_RNIHG744: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_ADD3\,
cout => N_58453,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_2\,
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_3_RNITN912: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIUCM01_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIV91B_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(6),
cin => N_58454);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_1_RNIRGA84: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_ADD3\,
cout => N_58455,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_3_RNIT8RT1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI1ULU_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIAP4A_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(32),
cin => N_58456);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_1_RNIMVN84: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_ADD3\,
cout => N_58457,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_3_RNI22152: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIPK9U_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIQDQB_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(31),
cin => N_58458);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_RNIPDME4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_ADD3\,
cout => N_58459,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_2_RNIDU962: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI8QA31_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIKUHA_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(30),
cin => N_58460);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_RNILEET4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_ADD3\,
cout => N_58461,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_3_RNI7CIF2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNID2U21_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIPLPE_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(29),
cin => N_58462);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_3_RNITV545: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_ADD3\,
cout => N_58463,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_2_RNIEURG2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIBC081_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIE80B_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(28),
cin => N_58464);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_2_RNI8LT55: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_ADD3\,
cout => N_58465,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_1_RNIE1MC2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIUEP31_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI8OUD_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(27),
cin => N_58466);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_3_RNID7VQ4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_ADD3\,
cout => N_58467,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_3_RNIDG992: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_2_RNI3RVV: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIDKIA_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(26),
cin => N_58468);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_2_RNIRDGB4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_ADD3\,
cout => N_58469,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_RNIB9RU1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI3LGT_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI0M77_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(25),
cin => N_58470);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_3_RNI09K04: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_ADD3\,
cout => N_58471,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_1_RNICBPP1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI8HOR_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIHCQB_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(24),
cin => N_58472);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_1_RNI90JT3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_ADD3\,
cout => N_58473,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_1_RNIH06V1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI3A9U_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIL8E8_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(23),
cin => N_58474);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_2_RNI2SU54: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_ADD3\,
cout => N_58475,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_3_RNIV6HT1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIFNFT_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI63Q6_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(22),
cin => N_58476);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_3_RNIP8L54: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_ADD3\,
cout => N_58477,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_RNI2D822: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIP4MS_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI8VDB_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(21),
cin => N_58478);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_2_RNIOKSC4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_ADD3\,
cout => N_58479,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_2_RNIQI402: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIB8E01_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIBR18_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(20),
cin => N_58480);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_3_RNI1EKR5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_ADD3\,
cout => N_58481,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_RNI1FN43: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIR65P1_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIJUEN_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(17),
cin => N_58482);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_1_RNIUTVU6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_ADD3\,
cout => N_58483,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_RNIDP8L3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_CARRY_1\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_2_RNI5GVM1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI532O_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(16),
cin => N_58484);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_3_RNIRECF7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_ADD3\,
cout => N_58485,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_RNIU49L3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNILRUS1_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIU9QO_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(15),
cin => N_58486);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_2_RNIGJC67: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_ADD3\,
cout => N_58487,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_1_RNI4U8C3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI31BD1_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNID8QB_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(14),
cin => N_58488);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_3_RNIFUB16: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_ADD3\,
cout => N_58489,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_RNITF8G2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI12SU_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIH4E8_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(13),
cin => N_58490);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_3_RNIKO8H4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_ADD3\,
cout => N_58491,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_RNIAO5S1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIH98P_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNICR88_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(12),
cin => N_58492);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_1_RNINFAL3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_ADD3\,
cout => N_58493,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_1_RNI37AK1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI9S2P_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIAN88_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(11),
cin => N_58494);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_3_RNITVDH3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_ADD3\,
cout => N_58495,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_RNIF89O1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIGV4R_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI6J88_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(10),
cin => N_58496);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_3_RNI0O5O3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_ADD3\,
cout => N_58497,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_RNI7V1R1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI2JRR_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI9M1B_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(9),
cin => N_58498);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_1_RNI31EU3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_ADD3\,
cout => N_58499,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_ADD2\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_V\(3),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_CARRY_2\);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_RNILHHU1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_ADD2\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_CARRY_2\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_ADD1\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_V\(2),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_CARRY_1\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIVHKU_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_ADD1\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_CARRY_1\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_ADD0\,
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_V\(1),
cin => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_CARRY_0\);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI6I1B_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_ADD0\,
cout => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_CARRY_0\,
dataa => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_V\(0),
datab => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.CTRLXERSHFT.SUMIN_5\(8),
cin => N_58500);
N_68349 <= not N_63;
N_68350 <= not \GRLFPC2_0.R.MK.BUSY_RET_5\;
N_68351 <= not \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_27_REP1: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO_REP1\,
d => N_58201,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_REP4_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP4\(0),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_REP3_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP3\(0),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_REP2_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(0),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_REP1_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(0),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_REP2_42_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(42),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_REP1_42_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(42),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_REP2_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP2\(15),
d => N_68351,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_REP1_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(15),
d => N_68351,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_REP2_17_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP2\(17),
d => N_58165,
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_REP1_17_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(17),
d => N_58165,
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_174: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(63),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(63),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_173: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(63),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(63),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_1: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN3_NOTXZYFROMD\,
d => N_58149,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_9: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN26_XZYBUSLSBS\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN26_XZYBUSLSBS_RETI\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_10: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5416\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.N_5416_RETI\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP0\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(15),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_15__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_171: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(62),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(62),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_170: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(62),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(62),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_168: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(61),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(61),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_167: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(61),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(61),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_165: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(64),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(64),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_164: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(64),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(64),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_162: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(77),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(77),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_161: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(77),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(77),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_159: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(69),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(69),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_158: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(69),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(69),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_156: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(68),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(68),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_155: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(68),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(68),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_153: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(67),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(67),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_152: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(67),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(67),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_150: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(76),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(76),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_149: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(76),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(76),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_147: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(75),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(75),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_146: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(75),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(75),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_145: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.FPI.LDOP_RETO\,
d => N_58150,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_144: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(74),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(74),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_143: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(74),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(74),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_141: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(73),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(73),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_140: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(73),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(73),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_138: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(72),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(72),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_137: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(72),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(72),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_135: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(71),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(71),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_134: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(71),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(71),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_69: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2_1\(9),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.EXPADDERSHFT.EXPYBUS_2_1_RETI\(9),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_REP1_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_REP1\(10),
d => N_58151,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_30_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(30),
d => N_58152,
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_133: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(8),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0_RETI\(8),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_8: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD\,
d => N_58153,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_7: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0\,
d => N_58154,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_48_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(48),
d => N_58155,
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_49_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(49),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(49),
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_132: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(7),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0_RETI\(7),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_50_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(50),
d => N_58156,
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_130: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_RETO\(70),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(70),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_129: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3_RETO\(70),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(70),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_128: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M14\(2),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M14_RETI\(2),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP0\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_104: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M14S2\,
d => N_58157,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP0\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_127: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_COUNTSUCCESSIVEZERO36_RETI\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP0\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_67: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WAITMULXFF.NOTSAMPLEDWAIT_RETO\,
d => N_58158,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_66: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_RETO\(4),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL\(4),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_10: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_PCTRL_NEW_1\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_126: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122\(4),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.DPATH_122_RETI\(4),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_53_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(53),
d => N_58159,
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_21_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(21),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(21),
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_125: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN8_TEMP_2\(0),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN8_TEMP_2_RETI\(0),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(1),
d => N_58160,
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_24_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(24),
d => N_58161,
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_124: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0\(5),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_0_RETI\(5),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_51_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(51),
d => N_58162,
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_52_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(52),
d => N_58163,
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_123: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS\(0),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS_RETI\(0),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RET_0: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.XZXBUS_2\(1),
d => N_58164,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(17),
d => N_58165,
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_115_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(115),
d => N_58166,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_122: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(16),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_RETI\(16),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_6: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD\,
d => N_58167,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_1: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN25_NOTXZYFROMD\,
d => N_58168,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_215_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(215),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(215),
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_121: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(15),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_RETI\(15),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_216_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(216),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(216),
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_120: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(14),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_RETI\(14),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_217_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(217),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(217),
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_119: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_13_M1_E\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_13_M1_E_RETI\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN15_NOTXZYFROMD_0_REP1\,
d => N_58169,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_16_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(16),
d => N_58170,
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_218_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(218),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(218),
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_118: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(12),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_RETI\(12),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_219_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(219),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(219),
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_117: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(11),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_RETI\(11),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_220_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(220),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(220),
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_116: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(10),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_RETI\(10),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_221_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(221),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(221),
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_115: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(9),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_RETI\(9),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_222_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(222),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(222),
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_114: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1\(8),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_RETI\(8),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_223_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(223),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(223),
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_113: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_3_M1_E_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_3_M1_E_1_RETI\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_228_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(228),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(228),
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_REP1_16_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_REP1\(16),
d => N_58171,
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_5_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(5),
d => N_58172,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_BUSY_RET: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => RST_RETO,
d => N_8,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_BUSY_RET_1: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.RST_RET_3\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.BUSYMULXFF.UN2_TEMP\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_64: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(79),
d => N_58173,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_0: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_62: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_RETO\(6),
d => N_58174,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_61: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.WQSTSETS_RETO\(4),
d => N_58175,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_60: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN14_CONDITIONAL_RETO\,
d => N_58176,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_58: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO(5),
d => N_62,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_2: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOINSTANDNOEXC_1\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_56: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO(6),
d => N_63,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_55: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_A13_7_1_RETO\(0),
d => N_58177,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_52: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO(9),
d => N_66,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_51: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_0_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN7_EXMIPTRLSBS_M_0\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_48: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO(12),
d => N_69,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_47: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(84),
d => N_58178,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_44: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO(11),
d => N_68,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_43: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_2_0_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTRESETORUNIMP_2_0\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_42: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28_RETO\,
d => N_58179,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_40: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO(8),
d => N_65,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_39: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_0_O19_2_RETO\(13),
d => N_58180,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_36: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO(10),
d => N_67,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_35: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M_0\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_112: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5\(1),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5_RETI\(1),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP0\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_13_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(13),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_13__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_11_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(11),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_11__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_12_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(12),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_12__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_111: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M2\(1),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M2_RETI\(1),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP0\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_17_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(17),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_17__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(15),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_15__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_16_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(16),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_16__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_110: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M8\(1),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M8_RETI\(1),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP0\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_9_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(9),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_9__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_7_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(7),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_7__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_8_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(8),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_8__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_109: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M11\(1),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M11_RETI\(1),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP0\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_5_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(5),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_5__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(3),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_3__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(4),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_4__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_108: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13_0\(3),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M13_0_RETI\(3),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP0\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_107: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12\(3),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M12_RETI\(3),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP0\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_26: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5S4\,
d => N_58181,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP0\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_23: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M11S4\,
d => N_58182,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP0\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(10),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_10__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_14_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(14),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_14__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_6_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(6),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M_0_6__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(2),
d => N_58183,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_100: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5\(0),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M5_RETI\(0),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP0\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_99: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M8\(0),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M8_RETI\(0),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP0\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_98: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M2\(0),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M2_RETI\(0),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP0\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_97: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M11\(0),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.COUNTSUCCESSIVEZERO_M11_RETI\(0),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN_REP0\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_96: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_6_M3_E\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_6_M3_E_RETI\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_RET: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN15_XZROUNDOUT\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN15_XZROUNDOUT_RETI\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_95: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM_A\(2),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_V_0_XX_MM_A_RETI\(2),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_2: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_REP1\,
d => N_58184,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_54_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(54),
d => N_58185,
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_94: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_372__G1_RETO\,
d => N_58186,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_91: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(113),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(113),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_89: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(85),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(85),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_20: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(85),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(85),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_86: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23_RETO\(84),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(84),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_21: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_REP1_RETO\,
d => N_58187,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_17: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(84),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(84),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_18: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_7_M3_E_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_7_M3_E_1_RETI\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_224_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(224),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(224),
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_225_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(225),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(225),
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_83: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_319__G1_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_319__G1\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_82: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.DPATH_NEW_7_SQMUXA_RETO\,
d => N_58188,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_81: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2_RETO\(60),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M2\(60),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_80: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_112__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_112__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_78: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_111__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_111__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_76: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_110__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_110__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_74: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_109__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_109__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_72: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_108__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_108__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_70: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_107__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_107__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_68: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_106__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_106__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_66: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_105__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_105__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_64: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_104__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_104__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_62: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_103__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_103__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_60: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_102__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_102__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_58: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_101__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_101__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_56: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_100__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_100__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_54: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_99__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_99__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_52: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_98__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_98__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_50: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_97__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_97__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_48: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_96__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_96__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_46: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_95__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_95__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_44: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_94__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_94__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_4: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_84__G0_I_A3_RETO\,
d => N_58189,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_43: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_93__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_93__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_42: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_92__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_92__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_41: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_91__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_91__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_40: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_90__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_90__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_39: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_89__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_89__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_38: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_88__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_88__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_37: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_87__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_87__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_35: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_86__G2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_0_86__G2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_33: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M4_0_RETI\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_0: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.UN16_NOTXZYFROMD_REP1\,
d => N_58190,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_32: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_4_M3_E\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_4_M3_E_RETI\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_31: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_SN_M2_RETI\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_5: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => RFO2_DATA1_RETO(27),
d => N_697,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_3: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => RFO2_DATA1_RETO(28),
d => N_698,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_16: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.EXTEND.TEMP_1\(1),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.EXTEND.TEMP_1_RETI\(1),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_8_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(8),
d => N_58191,
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_11_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(11),
d => N_58192,
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_58_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(58),
d => N_58193,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_25_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(25),
d => N_58194,
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_227_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(227),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(227),
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_RET_13: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_5_M3_E_1\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.FAX.TEMP_1_1_5_M3_E_1_RETI\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_226_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(226),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(226),
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_229_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(229),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(229),
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_55_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(55),
d => N_58195,
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_230_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(230),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(230),
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_56_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(56),
d => N_58196,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_57_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(57),
d => N_58197,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_231_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(231),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATHI\(231),
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_7: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP2\(0),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SUB_REP2_RETI\(0),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_19_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(19),
d => N_58198,
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_13_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(13),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(13),
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_9_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(9),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(9),
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_375_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(375),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_375__G0_0\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_72_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(72),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.NOTSQRTLFTCC_1_28\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_59_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(59),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_59__G0_XX_MM\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_29: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO\(2),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M\(2),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_23: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M_RETO\(4),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_I_M\(4),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_20: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_6_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_6\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_26: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_1_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_1\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_17: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_2_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_14: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_7_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_7\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_114_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(114),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_114__G0\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_83_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(83),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_X\(83),
clk => N_9,
clrn => VCC,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(83),
sload => \GRLFPC2_0.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_82_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(82),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_X\(82),
clk => N_9,
clrn => VCC,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(82),
sload => \GRLFPC2_0.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_81_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(81),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19_X\(81),
clk => N_9,
clrn => VCC,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(81),
sload => \GRLFPC2_0.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_80_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(80),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(80),
clk => N_9,
clrn => VCC,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(80),
sload => \GRLFPC2_0.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_79_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(79),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(79),
clk => N_9,
clrn => VCC,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(79),
sload => \GRLFPC2_0.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_78_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(78),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(78),
clk => N_9,
clrn => VCC,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(78),
sload => \GRLFPC2_0.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_66_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(66),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(66),
clk => N_9,
clrn => VCC,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(66),
sload => \GRLFPC2_0.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_65_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(65),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_19\(65),
clk => N_9,
clrn => VCC,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_M3\(65),
sload => \GRLFPC2_0.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_33: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_RETO\(6),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL\(6),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_32: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_C_RETO\,
d => N_58199,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_21: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_D_RETO\,
d => N_58200,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_30: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPI_D_INST_RETO(7),
d => N_64,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_28: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(54),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(54),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_27: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MULTIPLEXORMULXFF.UN10_SELECTEDMIPTR_RETO\,
d => N_58201,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_25: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_4_0_RETO\,
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_NOTSAMPLEDWAIT_1_4_0\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_22: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_U_RETO\(1),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_U\(1),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_19: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(53),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(53),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_16: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(0),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT\(0),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_12: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT_RETO\(3),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.RESULT\(3),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_8: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL_RETO\(3),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.PCTRL\(3),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_RET_4: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_RETO\(55),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(55),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_376_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(376),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_DIVMULTV\(0),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_12_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(12),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(12),
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_374_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(374),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_374__G0\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_14_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(14),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRLI\(14),
clk => N_9,
clrn => VCC,
ena => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_63_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(63),
d => \GRLFPC2_0.COMB.V.I.RES_1\(63),
clk => N_9,
clrn => VCC,
ena => G_8482,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_59_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(59),
d => \GRLFPC2_0.FPI.OP2_X\(62),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD7\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_58_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(58),
d => \GRLFPC2_0.FPI.OP2_X\(61),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD6\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_57_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(57),
d => \GRLFPC2_0.FPI.OP2_X\(60),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD5\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_56_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(56),
d => \GRLFPC2_0.FPI.OP2_X\(59),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD4\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_55_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(55),
d => \GRLFPC2_0.FPI.OP2_X\(58),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD3\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_54_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(54),
d => \GRLFPC2_0.FPI.OP2_X\(57),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD2\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_53_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(53),
d => \GRLFPC2_0.FPI.OP2_X\(56),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD1\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_52_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(52),
d => \GRLFPC2_0.FPI.OP2_X\(55),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD0\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_51_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(51),
d => \GRLFPC2_0.FPI.OP2_X\(54),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD54\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_50_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(50),
d => \GRLFPC2_0.FPI.OP2_X\(53),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD53\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_49_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(49),
d => \GRLFPC2_0.FPI.OP2_X\(52),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD52\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_48_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(48),
d => \GRLFPC2_0.FPI.OP2_X\(51),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD51\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_47_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(47),
d => \GRLFPC2_0.FPI.OP2_X\(50),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD50\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_46_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(46),
d => \GRLFPC2_0.FPI.OP2_X\(49),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD49\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_45_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(45),
d => \GRLFPC2_0.FPI.OP2_X\(48),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD48\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_44_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(44),
d => \GRLFPC2_0.FPI.OP2_X\(47),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD47\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_43_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(43),
d => \GRLFPC2_0.FPI.OP2_X\(46),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD46\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_42_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(42),
d => \GRLFPC2_0.FPI.OP2_X\(45),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD45\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_41_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(41),
d => \GRLFPC2_0.FPI.OP2_X\(44),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD44\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_40_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(40),
d => \GRLFPC2_0.FPI.OP2_X\(43),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD43\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_39_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(39),
d => \GRLFPC2_0.FPI.OP2_X\(42),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD42\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_38_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(38),
d => \GRLFPC2_0.FPI.OP2_X\(41),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD41\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_37_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(37),
d => \GRLFPC2_0.FPI.OP2_X\(40),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD40\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_36_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(36),
d => \GRLFPC2_0.FPI.OP2_X\(39),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD39\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_35_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(35),
d => \GRLFPC2_0.FPI.OP2_X\(38),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD38\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_34_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(34),
d => \GRLFPC2_0.FPI.OP2_X\(37),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD37\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_33_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(33),
d => \GRLFPC2_0.FPI.OP2_X\(36),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD36\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_32_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(32),
d => \GRLFPC2_0.FPI.OP2_X\(35),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD35\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_31_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(31),
d => \GRLFPC2_0.FPI.OP2_X\(34),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD34\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_30_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(30),
d => \GRLFPC2_0.FPI.OP2_X\(33),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD33\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_I_RES_29_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(29),
d => \GRLFPC2_0.FPI.OP2_X\(32),
clk => N_9,
clrn => VCC,
ena => G_8482,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD32\,
sload => \GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_116_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(116),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD57\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(118),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_117_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(117),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD56\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(119),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_118_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(118),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD55\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(120),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_119_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(119),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD54\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(121),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_120_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(120),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD53\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(122),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_121_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(121),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD52\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(123),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_122_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(122),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD51\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(124),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_123_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(123),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD50\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(125),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_124_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(124),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD49\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(126),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_125_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(125),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD48\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(127),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_126_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(126),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD47\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(128),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_127_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(127),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD46\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(129),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_128_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(128),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD45\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(130),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_129_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(129),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD44\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(131),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_130_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(130),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD43\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(132),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_131_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(131),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD42\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(133),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_132_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(132),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD41\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(134),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_133_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(133),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD40\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(135),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_134_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(134),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD39\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(136),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_135_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(135),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD38\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(137),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_136_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(136),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD37\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(138),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_137_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(137),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD36\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(139),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_138_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(138),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD35\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(140),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_139_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(139),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD34\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(141),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_140_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(140),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD33\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(142),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_141_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(141),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(141),
clk => N_9,
clrn => VCC,
ena => G_8368,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_142_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(142),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(142),
clk => N_9,
clrn => VCC,
ena => G_8368,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_143_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(143),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD30\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(145),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_144_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(144),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD29\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(146),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_145_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(145),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD28\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(147),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_146_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(146),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD27\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(148),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_147_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(147),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD26\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(149),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_148_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(148),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD25\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(150),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_149_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(149),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD24\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(151),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_150_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(150),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD23\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(152),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_151_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(151),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD22\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(153),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_152_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(152),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD21\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(154),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_153_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(153),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD20\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(155),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_154_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(154),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD19\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(156),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_155_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(155),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD18\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(157),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_156_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(156),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD17\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(158),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_157_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(157),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD16\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(159),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_158_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(158),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD15\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(160),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_159_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(159),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD14\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(161),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_160_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(160),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD13\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(162),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_161_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(161),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD12\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(163),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_162_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(162),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD11\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(164),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_163_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(163),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD10\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(165),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_164_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(164),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD9\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(166),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_165_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(165),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD8\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(167),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_166_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(166),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD7\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(168),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_167_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(167),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD6\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(169),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_168_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(168),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD5\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(170),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_169_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(169),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD4\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(171),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_170_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(170),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD3\,
clk => N_9,
clrn => VCC,
ena => G_8368,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(172),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_171_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(171),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(171),
clk => N_9,
clrn => VCC,
ena => G_8368,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_172_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(172),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(172),
clk => N_9,
clrn => VCC,
ena => G_8368,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_237_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(237),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_237__G0\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPAREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_238_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(238),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_238__G0\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPAREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_239_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(239),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_239__G0\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPAREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_240_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(240),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_240__G0\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPAREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_241_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(241),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_241__G0\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPAREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_242_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(242),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_242__G0\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPAREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_243_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(243),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_243__G0\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPAREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_244_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(244),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_244__G0\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPAREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_247_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(247),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(247),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_248_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(248),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(248),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_249_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(249),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(249),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_250_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(250),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(250),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_251_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(251),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(251),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_252_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(252),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(252),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_253_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(253),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(253),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_254_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(254),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(254),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_255_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(255),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(255),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_256_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(256),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(256),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_257_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(257),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(257),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_77_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(77),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW\(77),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_76_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(76),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_76__G0\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_74_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(74),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_0_0_74__G0\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_73_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(73),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.STARTSHFT.UN3_NOTRESETORUNIMP\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_71_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(71),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.UN36_PCTRL_NEW_I_0_G0\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_70_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(70),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(68),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_68_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(68),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.STARTSHFT.UN2_NOTDECODEDUNIMP\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_67_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(67),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.MAPMULXFF.UNIMPMAP_X\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW_6_0_67__G0_I_O4\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_66_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(66),
d => \GRLFPC2_0.FPI.START\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_65_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(65),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.PXS.PCTRL_NEW_2_0_65__G0\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_64_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(64),
d => N_58202,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_63_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(63),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_63__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_62_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(62),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_62__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_61_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(61),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_61__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_60_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(60),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_60__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_59_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(59),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_59__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_58_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(58),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_58__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_57_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(57),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_0_0\(56),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_56_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(56),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_56__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_55_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(55),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_55__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_54_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(54),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_54__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_53_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(53),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_53__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_52_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(52),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_52__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_51_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(51),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_51__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_50_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(50),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_50__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_49_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(49),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_49__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_48_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(48),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_19_0_I_I_I_0\(47),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_47_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(47),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_47__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_46_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(46),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_46__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_45_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(45),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_45__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_44_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(44),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_44__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_43_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(43),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_43__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_42_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(42),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_42__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_41_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(41),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_41__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_40_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(40),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_40__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_39_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(39),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_39__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_38_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(38),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_16_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(16),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_SCTRL_NEW_0_0__G0_I_M2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(15),
d => N_68351,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_14_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(14),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_I_0_0__G0\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_13_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(13),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_0_0_13__G0\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_12_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(12),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_R.SCTRL_2_IV\(0),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_11_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(11),
d => N_68349,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(10),
d => N_58203,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_9_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(9),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.UN17_U_RDN_I_0_8204_I_A2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_8_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(8),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.U_RDN_1_8221\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.RNDMODESELECT.TEMP\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_7_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(7),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW_0_0_7__G0\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(4),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW_0_0_7__G1\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(2),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_0_0_2__G0\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(1),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL_0_0_1__G0\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.SCTRL\(0),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.SXC.SCTRL_NEW_6_0_0__G0\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_36_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(36),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_36__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_35_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(35),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_35__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_34_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(34),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_34__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_33_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(33),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_33__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_32_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(32),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_32__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_31_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(31),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_31__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_29_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(29),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_29__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_28_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(28),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_28__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_27_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(27),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_27__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_26_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(26),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_26__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_25_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(25),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_25__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_24_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(24),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_24__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_23_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(23),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_23__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_22_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(22),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_22__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_21_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(21),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_21__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_20_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(20),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_20__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_18_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(18),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_18__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_7_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(7),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_7__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_6_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(6),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_6__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_5_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(5),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_5__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(4),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_4__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(3),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_3__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(2),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_2__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(1),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_1__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL\(0),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.PCTRL_2_0_0__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.PCTRL_NEW_21_0_38__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_377_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(377),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN1_GRFPUF_0\(0),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_373_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(373),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN2_MIXOIN_3\(0),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_372_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(372),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_372__G1\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_371_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(371),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(112),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_370_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(370),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(111),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_369_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(369),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(110),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_368_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(368),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(109),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_367_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(367),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(108),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_366_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(366),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(107),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_365_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(365),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(106),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_364_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(364),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(105),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_363_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(363),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(104),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_362_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(362),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(103),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_361_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(361),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(102),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_360_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(360),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(101),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_359_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(359),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(100),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_358_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(358),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(99),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP4\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_357_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(357),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(98),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_356_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(356),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(97),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_355_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(355),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(96),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_354_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(354),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(95),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_353_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(353),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(94),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_352_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(352),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(93),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_351_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(351),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(92),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_350_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(350),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(91),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_349_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(349),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(90),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_348_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(348),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(89),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_347_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(347),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(88),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_346_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(346),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(87),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_345_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(345),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(86),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_344_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(344),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(85),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_343_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(343),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(84),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_342_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(342),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(83),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_341_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(341),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(82),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_340_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(340),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(81),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_339_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(339),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(80),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_338_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(338),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(79),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_337_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(337),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(78),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_336_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(336),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(77),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_335_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(335),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(76),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_334_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(334),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(75),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_333_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(333),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(74),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_332_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(332),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(73),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_331_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(331),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(72),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP3\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_330_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(330),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(71),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_329_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(329),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(70),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_328_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(328),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(69),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_327_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(327),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(68),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_326_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(326),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(67),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_325_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(325),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(66),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_324_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(324),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(65),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_323_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(323),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(64),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_322_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(322),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(63),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_321_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(321),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(62),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_320_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(320),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_23\(61),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_319_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(319),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_319__G1\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_318_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(318),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_318__G1\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_317_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(317),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_317__G1\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_316_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(316),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_316__G1\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_315_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(315),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_315__G1\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_314_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(314),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_55_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_313_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(313),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_54_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_312_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(312),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_53_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_311_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(311),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_52_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_310_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(310),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_51_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_309_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(309),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_50_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_308_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(308),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_49_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_307_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(307),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_48_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_306_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(306),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_47_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_305_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(305),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_46_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_304_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(304),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_45_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP2\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_303_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(303),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_44_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_302_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(302),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_43_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_301_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(301),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_42_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_300_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(300),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_41_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_299_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(299),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_40_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_298_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(298),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_39_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_297_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(297),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_38_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_296_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(296),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_37_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_295_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(295),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_36_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_294_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(294),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_35_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_293_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(293),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_34_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_292_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(292),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_33_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_291_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(291),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_32_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_290_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(290),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_31_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_289_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(289),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_30_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_288_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(288),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_29_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_287_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(287),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_28_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_286_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(286),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_27_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_285_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(285),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_26_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_284_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(284),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_25_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_283_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(283),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_24_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_282_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(282),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_23_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_281_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(281),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_22_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_280_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(280),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_21_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_279_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(279),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_20_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_278_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(278),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_19_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_277_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(277),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_18_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB_REP1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_276_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(276),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_17_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_275_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(275),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_16_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_274_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(274),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_15_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_273_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(273),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_14_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_272_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(272),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_13_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_271_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(271),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_12_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_270_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(270),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_11_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_269_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(269),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_10_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_268_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(268),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_9_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_267_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(267),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_8_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_266_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(266),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_7_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_265_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(265),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_6_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_264_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(264),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_5_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_263_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(263),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.TRFWWRRAY.55.CI_4_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_262_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(262),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_262__G0_I_X4_0\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_261_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(261),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_261__G0_I_X4_0_0\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_260_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(260),
d => N_58204,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_259_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(259),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.DPATH_NEW_50_1.SUM_0\(0),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_258_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(258),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_258__G0_I_X4_0_0_0_1\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_246_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(246),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(246),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_245_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(245),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH\(245),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_236_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(236),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_236__G0\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_235_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(235),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_235__G0\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_234_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(234),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_234__G0\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_233_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(233),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_233__G0\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_232_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(232),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_3_232__G0\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_214_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(214),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD17\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_213_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(213),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD18\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_212_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(212),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD19\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_211_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(211),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD20\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_210_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(210),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD21\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_209_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(209),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD22\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_208_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(208),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD23\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_207_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(207),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD24\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_206_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(206),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD25\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_205_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(205),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD26\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_204_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(204),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD27\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_203_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(203),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD28\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_202_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(202),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD29\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_201_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(201),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD30\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_200_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(200),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD31\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_199_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(199),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD32\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_198_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(198),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD33\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_197_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(197),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD34\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_196_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(196),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD35\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_195_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(195),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD36\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_194_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(194),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD37\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_193_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(193),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD38\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_192_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(192),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD39\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_191_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(191),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD40\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_190_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(190),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD41\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_189_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(189),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD42\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_188_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(188),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD43\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_187_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(187),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD44\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_186_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(186),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD45\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_185_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(185),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD46\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_184_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(184),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD47\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_183_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(183),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD48\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_182_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(182),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD49\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_181_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(181),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD50\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_180_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(180),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD51\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_179_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(179),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD52\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_178_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(178),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD53\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_177_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(177),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD54\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_176_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(176),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD55\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_175_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(175),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD56\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_174_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(174),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD57\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_173_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(173),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_173__G0\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_47_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(47),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(47),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(47),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_46_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(46),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(46),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(46),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_45_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(45),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(45),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(45),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_44_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(44),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(44),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(44),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_43_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(43),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(43),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(43),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_42_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(42),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(42),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(42),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_41_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(41),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(41),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(41),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_40_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(40),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(40),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(40),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_39_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(39),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(39),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(39),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_38_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(38),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(38),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(38),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_37_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(37),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(37),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(37),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_36_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(36),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(36),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(36),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_35_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(35),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(35),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(35),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_34_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(34),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(34),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(34),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_33_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(33),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(33),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(33),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_32_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(32),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(32),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(32),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_31_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(31),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(31),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(31),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_30_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(30),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(30),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(30),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_29_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(29),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(29),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(29),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_28_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(28),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(28),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(28),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_27_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(27),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(27),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(27),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_26_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(26),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(26),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(26),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_23_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(23),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(23),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(23),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_22_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(22),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(22),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(22),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_20_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(20),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(20),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(20),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_19_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(19),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(19),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(19),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_18_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(18),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(18),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(18),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.R.DPATH\(0),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_4\(0),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_5\(0),
sload => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
GRLFPC2_0_R_MK_HOLDN2: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.HOLDN2\,
d => N_68350,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_LDOP_RET: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.LDOP_RET\,
d => N_17,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_LDOP_RET_3: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.LDOP_RET_3\,
d => N_58206,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_LDOP_RET_6: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.LDOP_RET_6\,
d => N_18,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_RST2: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.RST2\,
d => N_58207,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_RST_RET: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.RST_RET\,
d => N_58208,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_RST_RET_6: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.RST_RET_6\,
d => \GRLFPC2_0.R.MK.HOLDN2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_RST_RET_2: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.RST_RET_2\,
d => \GRLFPC2_0.R.MK.RST2\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_I_V: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.V\,
d => \GRLFPC2_0.R.I.V_1_0_G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.V_1_0_G0_I_O4\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_M_AFQ_RET_1: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.M.AFQ_RET_1\,
d => \GRLFPC2_0.COMB.UN1_FPCI_2_X\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_E_AFQ_RET_1: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.E.AFQ_RET_1\,
d => \GRLFPC2_0.COMB.UN3_HOLDN_X\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_M_AFQ_RET: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.M.AFQ_RET\,
d => \GRLFPC2_0.R.M.AFQ_RET_0_0_G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_M_AFSR_RET: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.M.AFSR_RET\,
d => \GRLFPC2_0.R.M.AFSR_RET_0_0_G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_A_RS2D: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RS2D\,
d => \GRLFPC2_0.R.A.RS2D_0_0_G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_A_RS1D: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RS1D\,
d => \GRLFPC2_0.COMB.RS1D_1_U\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_A_SEQERR_RET_3: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.SEQERR_RET_3\,
d => \GRLFPC2_0.N_1213_I_0_O2\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_M_SEQERR: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.M.SEQERR\,
d => \GRLFPC2_0.R.E.SEQERR\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_I_PC_RET_60: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_60\,
d => \GRLFPC2_0.R.I.RDD_0_0_G1_0_8238_I_O4\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_A_AFQ_RET_5: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.AFQ_RET_5\,
d => N_18,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_E_AFQ_RET: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.E.AFQ_RET\,
d => \GRLFPC2_0.COMB.V.A.AFQ_1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_A_ST_RET: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.ST_RET\,
d => \GRLFPC2_0.R.A.ST_RET_0_0_G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_E_SEQERR: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.E.SEQERR\,
d => \GRLFPC2_0.R.E.SEQERR_0_0_G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_E_AFSR_RET: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.E.AFSR_RET\,
d => \GRLFPC2_0.COMB.V.A.AFSR_1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_A_AFQ_RET_2: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.AFQ_RET_2\,
d => \GRLFPC2_0.N_939_I_I_A2\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_X_RDD: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.X.RDD\,
d => \GRLFPC2_0.R.M.RDD\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_M_RDD: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.M.RDD\,
d => \GRLFPC2_0.R.E.RDD\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_E_RDD: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.E.RDD\,
d => \GRLFPC2_0.R.A.RDD\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_A_RDD: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RDD\,
d => \GRLFPC2_0.R.A.RDD_0_0_G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_X_SEQERR: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.X.SEQERR\,
d => \GRLFPC2_0.R.M.SEQERR\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_A_LD: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.LD\,
d => \GRLFPC2_0.R.A.LD_0_0_G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_A_FPOP: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.FPOP\,
d => \GRLFPC2_0.R.A.FPOP_0_0_G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_I_EXEC: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.EXEC\,
d => \GRLFPC2_0.R.I.EXEC_0_0_G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_FTT_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.FTT\(2),
d => \GRLFPC2_0.R.FSR.FTT_0_0_2__G1_X\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_FTT_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.FTT\(0),
d => \GRLFPC2_0.R.FSR.FTT_0_0_0__G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_FSR_NONSTD: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.NONSTD\,
d => \GRLFPC2_0.R.FSR.NONSTD_0_0_G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_I_RDD: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RDD\,
d => \GRLFPC2_0.R.I.RDD_0_0_G1_0_8238_I\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_X_LD: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.X.LD\,
d => \GRLFPC2_0.R.X.LD_0_0_G1_X\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_X_FPOP: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.X.FPOP\,
d => \GRLFPC2_0.R.X.FPOP_0_0_G1_X\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_X_AFSR: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.X.AFSR\,
d => \GRLFPC2_0.R.X.AFSR_0_0_G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_X_AFQ: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.X.AFQ\,
d => \GRLFPC2_0.R.X.AFQ_0_0_G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_M_LD: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.M.LD\,
d => \GRLFPC2_0.R.M.LD_0_0_G1_X\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_M_FPOP: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.M.FPOP\,
d => \GRLFPC2_0.R.M.FPOP_0_0_G1_X\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_E_LD: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.E.LD\,
d => \GRLFPC2_0.R.E.LD_0_0_G1_X\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_E_FPOP: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.E.FPOP\,
d => \GRLFPC2_0.R.E.FPOP_0_0_G1_X\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_BUSY2_RET: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.BUSY2_RET\,
d => \GRLFPC2_0.R.MK.BUSY2_RET_0_0_A2_0_G0_X\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_BUSY_RET_3: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.BUSY_RET_3\,
d => \GRLFPC2_0.R.MK.BUSY_RET_3_0_0_A2_X\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_BUSY_RET_2: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.BUSY_RET_2\,
d => \GRLFPC2_0.R.MK.BUSY_RET_2_0_0_A2_0_G0_X\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_BUSY2_RET_1: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.BUSY2_RET_1\,
d => \GRLFPC2_0.R.MK.BUSY2_RET_1_0_0_A2_0_G0\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_BUSY_RET_5: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.BUSY_RET_5\,
d => \GRLFPC2_0.R.MK.HOLDN1_0_I_A2_X\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC2_0_R_MK_BUSY_RET_4: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.BUSY_RET_4\,
d => \GRLFPC2_0.R.MK.BUSY_RET_4_0_0_A2_0_G0\,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(0),
d => N_333,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(1),
d => N_334,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(2),
d => N_335,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(3),
d => N_336,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(4),
d => N_337,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_5_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(5),
d => N_338,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_6_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(6),
d => N_339,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_7_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(7),
d => N_340,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_8_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(8),
d => N_341,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_9_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(9),
d => N_342,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(10),
d => N_343,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_11_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(11),
d => N_344,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_12_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(12),
d => N_345,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_13_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(13),
d => N_346,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_14_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(14),
d => N_347,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(15),
d => N_348,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_16_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(16),
d => N_349,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_17_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(17),
d => N_350,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_18_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(18),
d => N_351,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_19_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(19),
d => N_352,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_20_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(20),
d => N_353,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_21_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(21),
d => N_354,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_22_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(22),
d => N_355,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_23_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(23),
d => N_356,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_24_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(24),
d => N_357,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_25_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(25),
d => N_358,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_26_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(26),
d => N_359,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_27_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(27),
d => N_360,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_28_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(28),
d => N_361,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_29_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(29),
d => N_362,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_30_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(30),
d => N_363,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_INST_31_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.INST\(31),
d => N_364,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.INST_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_E_STDATA_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(0),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(0),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(0),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(1),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(1),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(1),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(2),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(2),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(2),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(3),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(3),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(3),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(4),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(4),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(4),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_5_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(5),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(5),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(5),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_6_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(6),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(6),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(6),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_7_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(7),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(7),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(7),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_8_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(8),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(8),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(8),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_9_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(9),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(9),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(9),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(10),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(10),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(10),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_11_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(11),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(11),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(11),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_12_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(12),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(12),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(12),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_13_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(13),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(13),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(13),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_14_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(14),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(14),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(14),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(15),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(15),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(15),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_16_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(16),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(16),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(16),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_17_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(17),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(17),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(17),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_18_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(18),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(18),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(18),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_19_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(19),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(19),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(19),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_20_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(20),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(20),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(20),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_21_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(21),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(21),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(21),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_22_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(22),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(22),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(22),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_23_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(23),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(23),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(23),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_24_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(24),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(24),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(24),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_25_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(25),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(25),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(25),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_26_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(26),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(26),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(26),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_27_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(27),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(27),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(27),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_28_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(28),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(28),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(28),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_29_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(29),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(29),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(29),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_30_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(30),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(30),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(30),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_E_STDATA_31_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_DATAZ(31),
d => \GRLFPC2_0.COMB.V.E.STDATA_1_0_X\(31),
clk => N_9,
clrn => VCC,
ena => N_17,
asdata => \GRLFPC2_0.COMB.V.E.STDATA_1_1\(31),
sload => \GRLFPC2_0.COMB.V.A.AFQ_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC2_0_R_FSR_RD_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.RD\(0),
d => \GRLFPC2_0.R.FSR.RD_0_0_0__G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_RD_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.RD\(1),
d => \GRLFPC2_0.R.FSR.RD_0_0_1__G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_TEM_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.TEM\(0),
d => \GRLFPC2_0.R.FSR.TEM_1_0_0__G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_TEM_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.TEM\(1),
d => \GRLFPC2_0.R.FSR.TEM_1_0_1__G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_TEM_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.TEM\(2),
d => \GRLFPC2_0.R.FSR.TEM_1_0_2__G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_TEM_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.TEM\(3),
d => \GRLFPC2_0.R.FSR.TEM_1_0_3__G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_TEM_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.TEM\(4),
d => \GRLFPC2_0.R.FSR.TEM_1_0_4__G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_STATE_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.STATE\(0),
d => \GRLFPC2_0.R.STATE_0_0_0__G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_STATE_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.STATE\(1),
d => \GRLFPC2_0.COMB.V.STATE_1_IV\(1),
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RF1REN_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RF1REN\(2),
d => \GRLFPC2_0.COMB.RF1REN_1_0_0\(2),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RF1REN_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RF1REN\(1),
d => \GRLFPC2_0.COMB.V.A.RF1REN_1_8259_I\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RF2REN_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RF2REN\(2),
d => \GRLFPC2_0.COMB.V.A.RF2REN_1_0_8287_I\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RF2REN_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RF2REN\(1),
d => \GRLFPC2_0.COMB.V.A.RF2REN_1_8311_I\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_FCC_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_CCZ(0),
d => \GRLFPC2_0.R.FSR.FCC_0_0_0__G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_FCC_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => CPO_CCZ(1),
d => \GRLFPC2_0.R.FSR.FCC_0_0_1__G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_AEXC_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.AEXC\(0),
d => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV\(0),
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_AEXC_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.AEXC\(1),
d => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV\(1),
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_AEXC_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.AEXC\(2),
d => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV\(2),
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_AEXC_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.AEXC\(3),
d => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV\(3),
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_AEXC_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.AEXC\(4),
d => \GRLFPC2_0.COMB.V.FSR.AEXC_1_IV\(4),
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_CEXC_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.CEXC\(0),
d => \GRLFPC2_0.R.FSR.CEXC_1_0_0__G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_CEXC_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.CEXC\(1),
d => \GRLFPC2_0.R.FSR.CEXC_1_0_1__G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_CEXC_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.CEXC\(2),
d => \GRLFPC2_0.R.FSR.CEXC_1_0_2__G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_CEXC_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.CEXC\(3),
d => \GRLFPC2_0.R.FSR.CEXC_1_0_3__G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_FSR_CEXC_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.FSR.CEXC\(4),
d => \GRLFPC2_0.R.FSR.CEXC_1_0_4__G1\,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_MOV_RET_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.MOV_RET\(0),
d => N_87,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_MOV_RET_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.MOV_RET\(2),
d => N_62,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_MOV_RET_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.MOV_RET\(3),
d => N_63,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_MOV_RET_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.MOV_RET\(4),
d => N_64,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_MOV_RET_5_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.MOV_RET\(5),
d => N_65,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_MOV_RET_6_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.MOV_RET\(6),
d => N_66,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_MOV_RET_7_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.MOV_RET\(7),
d => N_67,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_MOV_RET_8_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.MOV_RET\(8),
d => N_68,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_MOV_RET_9_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.MOV_RET\(9),
d => N_69,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_MOV_RET_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.MOV_RET\(10),
d => N_70,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_MOV_RET_11_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.MOV_RET\(11),
d => N_76,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_MOV_RET_12_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.MOV_RET\(12),
d => N_77,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_MOV_RET_13_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.MOV_RET\(13),
d => N_78,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_MOV_RET_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.MOV_RET\(15),
d => N_80,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_SEQERR_RET_4_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.SEQERR_RET_4\(0),
d => \GRLFPC2_0.R.STATE\(0),
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_SEQERR_RET_4_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.SEQERR_RET_4\(1),
d => \GRLFPC2_0.R.STATE\(1),
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_ST_RET_2_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.ST_RET_2\(0),
d => N_91,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_ST_RET_2_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.ST_RET_2\(1),
d => N_92,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_AFQ_RET_5_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.AFQ_RET\(5),
d => N_79,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_AFQ_RET_7_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.AFQ_RET\(7),
d => N_81,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_AFQ_RET_9_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.AFQ_RET\(9),
d => N_88,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_CC_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.CC\(0),
d => \GRLFPC2_0.R.I.CC_0_0_0__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_CC_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.CC\(1),
d => \GRLFPC2_0.R.I.CC_0_0_1__G2\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(0),
d => \GRLFPC2_0.R.I.PC_RET_30\(0),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(1),
d => \GRLFPC2_0.R.I.PC_RET_30\(1),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(2),
d => \GRLFPC2_0.R.I.PC_RET_30\(2),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(3),
d => \GRLFPC2_0.R.I.PC_RET_30\(3),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(4),
d => \GRLFPC2_0.R.I.PC_RET_30\(4),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_5_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(5),
d => \GRLFPC2_0.R.I.PC_RET_30\(5),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_6_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(6),
d => \GRLFPC2_0.R.I.PC_RET_30\(6),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_7_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(7),
d => \GRLFPC2_0.R.I.PC_RET_30\(7),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_8_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(8),
d => \GRLFPC2_0.R.I.PC_RET_30\(8),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_9_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(9),
d => \GRLFPC2_0.R.I.PC_RET_30\(9),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(10),
d => \GRLFPC2_0.R.I.PC_RET_30\(10),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_11_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(11),
d => \GRLFPC2_0.R.I.PC_RET_30\(11),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_12_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(12),
d => \GRLFPC2_0.R.I.PC_RET_30\(12),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_13_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(13),
d => \GRLFPC2_0.R.I.PC_RET_30\(13),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_14_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(14),
d => \GRLFPC2_0.R.I.PC_RET_30\(14),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(15),
d => \GRLFPC2_0.R.I.PC_RET_30\(15),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_16_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(16),
d => \GRLFPC2_0.R.I.PC_RET_30\(16),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_17_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(17),
d => \GRLFPC2_0.R.I.PC_RET_30\(17),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_18_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(18),
d => \GRLFPC2_0.R.I.PC_RET_30\(18),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_19_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(19),
d => \GRLFPC2_0.R.I.PC_RET_30\(19),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_20_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(20),
d => \GRLFPC2_0.R.I.PC_RET_30\(20),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_21_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(21),
d => \GRLFPC2_0.R.I.PC_RET_30\(21),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_22_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(22),
d => \GRLFPC2_0.R.I.PC_RET_30\(22),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_23_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(23),
d => \GRLFPC2_0.R.I.PC_RET_30\(23),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_24_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(24),
d => \GRLFPC2_0.R.I.PC_RET_30\(24),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_25_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(25),
d => \GRLFPC2_0.R.I.PC_RET_30\(25),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_26_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(26),
d => \GRLFPC2_0.R.I.PC_RET_30\(26),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_27_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(27),
d => \GRLFPC2_0.R.I.PC_RET_30\(27),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_28_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(28),
d => \GRLFPC2_0.R.I.PC_RET_30\(28),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_29_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET\(29),
d => \GRLFPC2_0.R.I.PC_RET_30\(29),
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.R.I.PC_RET_1_0_0__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(0),
d => N_303,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(1),
d => N_304,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(2),
d => N_305,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(3),
d => N_306,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(4),
d => N_307,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_5_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(5),
d => N_308,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_6_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(6),
d => N_309,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_7_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(7),
d => N_310,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_8_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(8),
d => N_311,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_9_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(9),
d => N_312,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(10),
d => N_313,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_11_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(11),
d => N_314,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_12_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(12),
d => N_315,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_13_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(13),
d => N_316,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_14_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(14),
d => N_317,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(15),
d => N_318,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_16_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(16),
d => N_319,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_17_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(17),
d => N_320,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_18_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(18),
d => N_321,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_19_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(19),
d => N_322,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_20_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(20),
d => N_323,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_21_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(21),
d => N_324,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_22_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(22),
d => N_325,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_23_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(23),
d => N_326,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_24_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(24),
d => N_327,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_25_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(25),
d => N_328,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_26_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(26),
d => N_329,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_27_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(27),
d => N_330,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_28_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(28),
d => N_331,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_PC_RET_30_29_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.PC_RET_30\(29),
d => N_332,
clk => N_9,
clrn => VCC,
ena => N_17,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_EXC_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.EXC\(0),
d => \GRLFPC2_0.R.I.EXC_0\(0),
clk => N_9,
clrn => VCC,
ena => G_8482,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_EXC_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.EXC\(1),
d => \GRLFPC2_0.R.I.EXC_2_0_1__G2\,
clk => N_9,
clrn => VCC,
ena => G_8482,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_EXC_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.EXC\(2),
d => \GRLFPC2_0.R.I.EXC_2_0_2__G2\,
clk => N_9,
clrn => VCC,
ena => G_8482,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_EXC_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.EXC\(3),
d => \GRLFPC2_0.R.I.EXC_2_0_3__G2\,
clk => N_9,
clrn => VCC,
ena => G_8482,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_EXC_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.EXC\(4),
d => \GRLFPC2_0.R.I.EXC_2_0_4__G2\,
clk => N_9,
clrn => VCC,
ena => G_8482,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_MK_LDOP_RET_4_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.LDOP_RET_4\(0),
d => \GRLFPC2_0.R.STATE\(0),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_MK_LDOP_RET_4_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.LDOP_RET_4\(1),
d => \GRLFPC2_0.R.STATE\(1),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_MK_LDOP_RET_1_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.LDOP_RET_1\(0),
d => N_91,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_MK_LDOP_RET_1_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.LDOP_RET_1\(1),
d => N_92,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_MK_LDOP_RET_1_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.LDOP_RET_1\(2),
d => N_81,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_MK_LDOP_RET_1_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.LDOP_RET_1\(3),
d => N_80,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_MK_LDOP_RET_1_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.LDOP_RET_1\(4),
d => N_79,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_MK_LDOP_RET_1_5_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.LDOP_RET_1\(5),
d => N_78,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_MK_LDOP_RET_1_6_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.LDOP_RET_1\(6),
d => N_77,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_MK_LDOP_RET_1_7_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.LDOP_RET_1\(7),
d => N_87,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_MK_LDOP_RET_1_8_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.MK.LDOP_RET_1\(8),
d => N_88,
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RS1_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RS1\(0),
d => \GRLFPC2_0.COMB.RS1_1\(0),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RS1_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RS1\(1),
d => \GRLFPC2_0.COMB.RS1_1\(1),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RS1_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RS1\(2),
d => \GRLFPC2_0.COMB.RS1_1\(2),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RS1_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RS1\(3),
d => \GRLFPC2_0.COMB.RS1_1\(3),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RS1_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RS1\(4),
d => \GRLFPC2_0.COMB.RS1_1\(4),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(0),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD3\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(1),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD4\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(2),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD5\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(3),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD6\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(4),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD7\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_5_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(5),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD8\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_6_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(6),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD9\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_7_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(7),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD10\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_8_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(8),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD11\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_9_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(9),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD12\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_10_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(10),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD13\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_11_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(11),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD14\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_12_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(12),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD15\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_13_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(13),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD16\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_14_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(14),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD17\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_15_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(15),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD18\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_16_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(16),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD19\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_17_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(17),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD20\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_18_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(18),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD21\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_19_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(19),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD22\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_20_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(20),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD23\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_21_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(21),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD24\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_22_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(22),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD25\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_23_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(23),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD26\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_24_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(24),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD27\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_25_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(25),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD28\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_26_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(26),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD29\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_27_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(27),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD30\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_28_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(28),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUF_ADD31\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_60_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(60),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD8\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_61_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(61),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD9\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_I_RES_62_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.I.RES\(62),
d => \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.UN6_GRFPUE_ADD10\,
clk => N_9,
clrn => VCC,
ena => \GRLFPC2_0.COMB.UN6_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RS2_0_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RS2\(0),
d => \GRLFPC2_0.COMB.RS2_1\(0),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RS2_1_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RS2\(1),
d => \GRLFPC2_0.COMB.RS2_1\(1),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RS2_2_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RS2\(2),
d => \GRLFPC2_0.COMB.RS2_1\(2),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RS2_3_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RS2\(3),
d => \GRLFPC2_0.COMB.RS2_1\(3),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC2_0_R_A_RS2_4_\: dffeas generic map (
    is_wysiwyg => "true")
port map (
q => \GRLFPC2_0.R.A.RS2\(4),
d => \GRLFPC2_0.COMB.RS2_1\(4),
clk => N_9,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
N_8 <= RST_INTERNAL;
N_9 <= CLK_INTERNAL;
N_17 <= HOLDN_INTERNAL;
N_18 <= CPI_FLUSH_INTERNAL;
N_19 <= CPI_EXACK_INTERNAL;
N_20 <= CPI_A_RS1_INTERNAL;
N_21 <= CPI_A_RS1_INTERNAL_0;
N_22 <= CPI_A_RS1_INTERNAL_1;
N_23 <= CPI_A_RS1_INTERNAL_2;
N_24 <= CPI_A_RS1_INTERNAL_3;
N_25 <= CPI_D_PC_INTERNAL;
N_26 <= CPI_D_PC_INTERNAL_0;
N_27 <= CPI_D_PC_INTERNAL_1;
N_28 <= CPI_D_PC_INTERNAL_2;
N_29 <= CPI_D_PC_INTERNAL_3;
N_30 <= CPI_D_PC_INTERNAL_4;
N_31 <= CPI_D_PC_INTERNAL_5;
N_32 <= CPI_D_PC_INTERNAL_6;
N_33 <= CPI_D_PC_INTERNAL_7;
N_34 <= CPI_D_PC_INTERNAL_8;
N_35 <= CPI_D_PC_INTERNAL_9;
N_36 <= CPI_D_PC_INTERNAL_10;
N_37 <= CPI_D_PC_INTERNAL_11;
N_38 <= CPI_D_PC_INTERNAL_12;
N_39 <= CPI_D_PC_INTERNAL_13;
N_40 <= CPI_D_PC_INTERNAL_14;
N_41 <= CPI_D_PC_INTERNAL_15;
N_42 <= CPI_D_PC_INTERNAL_16;
N_43 <= CPI_D_PC_INTERNAL_17;
N_44 <= CPI_D_PC_INTERNAL_18;
N_45 <= CPI_D_PC_INTERNAL_19;
N_46 <= CPI_D_PC_INTERNAL_20;
N_47 <= CPI_D_PC_INTERNAL_21;
N_48 <= CPI_D_PC_INTERNAL_22;
N_49 <= CPI_D_PC_INTERNAL_23;
N_50 <= CPI_D_PC_INTERNAL_24;
N_51 <= CPI_D_PC_INTERNAL_25;
N_52 <= CPI_D_PC_INTERNAL_26;
N_53 <= CPI_D_PC_INTERNAL_27;
N_54 <= CPI_D_PC_INTERNAL_28;
N_55 <= CPI_D_PC_INTERNAL_29;
N_56 <= CPI_D_PC_INTERNAL_30;
N_57 <= CPI_D_INST_INTERNAL;
N_58 <= CPI_D_INST_INTERNAL_0;
N_59 <= CPI_D_INST_INTERNAL_1;
N_60 <= CPI_D_INST_INTERNAL_2;
N_61 <= CPI_D_INST_INTERNAL_3;
N_62 <= CPI_D_INST_INTERNAL_4;
N_63 <= CPI_D_INST_INTERNAL_5;
N_64 <= CPI_D_INST_INTERNAL_6;
N_65 <= CPI_D_INST_INTERNAL_7;
N_66 <= CPI_D_INST_INTERNAL_8;
N_67 <= CPI_D_INST_INTERNAL_9;
N_68 <= CPI_D_INST_INTERNAL_10;
N_69 <= CPI_D_INST_INTERNAL_11;
N_70 <= CPI_D_INST_INTERNAL_12;
N_71 <= CPI_D_INST_INTERNAL_13;
N_72 <= CPI_D_INST_INTERNAL_14;
N_73 <= CPI_D_INST_INTERNAL_15;
N_74 <= CPI_D_INST_INTERNAL_16;
N_75 <= CPI_D_INST_INTERNAL_17;
N_76 <= CPI_D_INST_INTERNAL_18;
N_77 <= CPI_D_INST_INTERNAL_19;
N_78 <= CPI_D_INST_INTERNAL_20;
N_79 <= CPI_D_INST_INTERNAL_21;
N_80 <= CPI_D_INST_INTERNAL_22;
N_81 <= CPI_D_INST_INTERNAL_23;
N_82 <= CPI_D_INST_INTERNAL_24;
N_83 <= CPI_D_INST_INTERNAL_25;
N_84 <= CPI_D_INST_INTERNAL_26;
N_85 <= CPI_D_INST_INTERNAL_27;
N_86 <= CPI_D_INST_INTERNAL_28;
N_87 <= CPI_D_INST_INTERNAL_29;
N_88 <= CPI_D_INST_INTERNAL_30;
N_89 <= CPI_D_CNT_INTERNAL;
N_90 <= CPI_D_CNT_INTERNAL_0;
N_91 <= CPI_D_TRAP_INTERNAL;
N_92 <= CPI_D_ANNUL_INTERNAL;
N_93 <= CPI_D_PV_INTERNAL;
N_94 <= CPI_A_PC_INTERNAL;
N_95 <= CPI_A_PC_INTERNAL_0;
N_96 <= CPI_A_PC_INTERNAL_1;
N_97 <= CPI_A_PC_INTERNAL_2;
N_98 <= CPI_A_PC_INTERNAL_3;
N_99 <= CPI_A_PC_INTERNAL_4;
N_100 <= CPI_A_PC_INTERNAL_5;
N_101 <= CPI_A_PC_INTERNAL_6;
N_102 <= CPI_A_PC_INTERNAL_7;
N_103 <= CPI_A_PC_INTERNAL_8;
N_104 <= CPI_A_PC_INTERNAL_9;
N_105 <= CPI_A_PC_INTERNAL_10;
N_106 <= CPI_A_PC_INTERNAL_11;
N_107 <= CPI_A_PC_INTERNAL_12;
N_108 <= CPI_A_PC_INTERNAL_13;
N_109 <= CPI_A_PC_INTERNAL_14;
N_110 <= CPI_A_PC_INTERNAL_15;
N_111 <= CPI_A_PC_INTERNAL_16;
N_112 <= CPI_A_PC_INTERNAL_17;
N_113 <= CPI_A_PC_INTERNAL_18;
N_114 <= CPI_A_PC_INTERNAL_19;
N_115 <= CPI_A_PC_INTERNAL_20;
N_116 <= CPI_A_PC_INTERNAL_21;
N_117 <= CPI_A_PC_INTERNAL_22;
N_118 <= CPI_A_PC_INTERNAL_23;
N_119 <= CPI_A_PC_INTERNAL_24;
N_120 <= CPI_A_PC_INTERNAL_25;
N_121 <= CPI_A_PC_INTERNAL_26;
N_122 <= CPI_A_PC_INTERNAL_27;
N_123 <= CPI_A_PC_INTERNAL_28;
N_124 <= CPI_A_PC_INTERNAL_29;
N_125 <= CPI_A_PC_INTERNAL_30;
N_126 <= CPI_A_INST_INTERNAL;
N_127 <= CPI_A_INST_INTERNAL_0;
N_128 <= CPI_A_INST_INTERNAL_1;
N_129 <= CPI_A_INST_INTERNAL_2;
N_130 <= CPI_A_INST_INTERNAL_3;
N_131 <= CPI_A_INST_INTERNAL_4;
N_132 <= CPI_A_INST_INTERNAL_5;
N_133 <= CPI_A_INST_INTERNAL_6;
N_134 <= CPI_A_INST_INTERNAL_7;
N_135 <= CPI_A_INST_INTERNAL_8;
N_136 <= CPI_A_INST_INTERNAL_9;
N_137 <= CPI_A_INST_INTERNAL_10;
N_138 <= CPI_A_INST_INTERNAL_11;
N_139 <= CPI_A_INST_INTERNAL_12;
N_140 <= CPI_A_INST_INTERNAL_13;
N_141 <= CPI_A_INST_INTERNAL_14;
N_142 <= CPI_A_INST_INTERNAL_15;
N_143 <= CPI_A_INST_INTERNAL_16;
N_144 <= CPI_A_INST_INTERNAL_17;
N_145 <= CPI_A_INST_INTERNAL_18;
N_146 <= CPI_A_INST_INTERNAL_19;
N_147 <= CPI_A_INST_INTERNAL_20;
N_148 <= CPI_A_INST_INTERNAL_21;
N_149 <= CPI_A_INST_INTERNAL_22;
N_150 <= CPI_A_INST_INTERNAL_23;
N_151 <= CPI_A_INST_INTERNAL_24;
N_152 <= CPI_A_INST_INTERNAL_25;
N_153 <= CPI_A_INST_INTERNAL_26;
N_154 <= CPI_A_INST_INTERNAL_27;
N_155 <= CPI_A_INST_INTERNAL_28;
N_156 <= CPI_A_INST_INTERNAL_29;
N_157 <= CPI_A_INST_INTERNAL_30;
N_158 <= CPI_A_CNT_INTERNAL;
N_159 <= CPI_A_CNT_INTERNAL_0;
N_160 <= CPI_A_TRAP_INTERNAL;
N_161 <= CPI_A_ANNUL_INTERNAL;
N_162 <= CPI_A_PV_INTERNAL;
N_163 <= CPI_E_PC_INTERNAL;
N_164 <= CPI_E_PC_INTERNAL_0;
N_165 <= CPI_E_PC_INTERNAL_1;
N_166 <= CPI_E_PC_INTERNAL_2;
N_167 <= CPI_E_PC_INTERNAL_3;
N_168 <= CPI_E_PC_INTERNAL_4;
N_169 <= CPI_E_PC_INTERNAL_5;
N_170 <= CPI_E_PC_INTERNAL_6;
N_171 <= CPI_E_PC_INTERNAL_7;
N_172 <= CPI_E_PC_INTERNAL_8;
N_173 <= CPI_E_PC_INTERNAL_9;
N_174 <= CPI_E_PC_INTERNAL_10;
N_175 <= CPI_E_PC_INTERNAL_11;
N_176 <= CPI_E_PC_INTERNAL_12;
N_177 <= CPI_E_PC_INTERNAL_13;
N_178 <= CPI_E_PC_INTERNAL_14;
N_179 <= CPI_E_PC_INTERNAL_15;
N_180 <= CPI_E_PC_INTERNAL_16;
N_181 <= CPI_E_PC_INTERNAL_17;
N_182 <= CPI_E_PC_INTERNAL_18;
N_183 <= CPI_E_PC_INTERNAL_19;
N_184 <= CPI_E_PC_INTERNAL_20;
N_185 <= CPI_E_PC_INTERNAL_21;
N_186 <= CPI_E_PC_INTERNAL_22;
N_187 <= CPI_E_PC_INTERNAL_23;
N_188 <= CPI_E_PC_INTERNAL_24;
N_189 <= CPI_E_PC_INTERNAL_25;
N_190 <= CPI_E_PC_INTERNAL_26;
N_191 <= CPI_E_PC_INTERNAL_27;
N_192 <= CPI_E_PC_INTERNAL_28;
N_193 <= CPI_E_PC_INTERNAL_29;
N_194 <= CPI_E_PC_INTERNAL_30;
N_195 <= CPI_E_INST_INTERNAL;
N_196 <= CPI_E_INST_INTERNAL_0;
N_197 <= CPI_E_INST_INTERNAL_1;
N_198 <= CPI_E_INST_INTERNAL_2;
N_199 <= CPI_E_INST_INTERNAL_3;
N_200 <= CPI_E_INST_INTERNAL_4;
N_201 <= CPI_E_INST_INTERNAL_5;
N_202 <= CPI_E_INST_INTERNAL_6;
N_203 <= CPI_E_INST_INTERNAL_7;
N_204 <= CPI_E_INST_INTERNAL_8;
N_205 <= CPI_E_INST_INTERNAL_9;
N_206 <= CPI_E_INST_INTERNAL_10;
N_207 <= CPI_E_INST_INTERNAL_11;
N_208 <= CPI_E_INST_INTERNAL_12;
N_209 <= CPI_E_INST_INTERNAL_13;
N_210 <= CPI_E_INST_INTERNAL_14;
N_211 <= CPI_E_INST_INTERNAL_15;
N_212 <= CPI_E_INST_INTERNAL_16;
N_213 <= CPI_E_INST_INTERNAL_17;
N_214 <= CPI_E_INST_INTERNAL_18;
N_215 <= CPI_E_INST_INTERNAL_19;
N_216 <= CPI_E_INST_INTERNAL_20;
N_217 <= CPI_E_INST_INTERNAL_21;
N_218 <= CPI_E_INST_INTERNAL_22;
N_219 <= CPI_E_INST_INTERNAL_23;
N_220 <= CPI_E_INST_INTERNAL_24;
N_221 <= CPI_E_INST_INTERNAL_25;
N_222 <= CPI_E_INST_INTERNAL_26;
N_223 <= CPI_E_INST_INTERNAL_27;
N_224 <= CPI_E_INST_INTERNAL_28;
N_225 <= CPI_E_INST_INTERNAL_29;
N_226 <= CPI_E_INST_INTERNAL_30;
N_227 <= CPI_E_CNT_INTERNAL;
N_228 <= CPI_E_CNT_INTERNAL_0;
N_229 <= CPI_E_TRAP_INTERNAL;
N_230 <= CPI_E_ANNUL_INTERNAL;
N_231 <= CPI_E_PV_INTERNAL;
N_232 <= CPI_M_PC_INTERNAL;
N_233 <= CPI_M_PC_INTERNAL_0;
N_234 <= CPI_M_PC_INTERNAL_1;
N_235 <= CPI_M_PC_INTERNAL_2;
N_236 <= CPI_M_PC_INTERNAL_3;
N_237 <= CPI_M_PC_INTERNAL_4;
N_238 <= CPI_M_PC_INTERNAL_5;
N_239 <= CPI_M_PC_INTERNAL_6;
N_240 <= CPI_M_PC_INTERNAL_7;
N_241 <= CPI_M_PC_INTERNAL_8;
N_242 <= CPI_M_PC_INTERNAL_9;
N_243 <= CPI_M_PC_INTERNAL_10;
N_244 <= CPI_M_PC_INTERNAL_11;
N_245 <= CPI_M_PC_INTERNAL_12;
N_246 <= CPI_M_PC_INTERNAL_13;
N_247 <= CPI_M_PC_INTERNAL_14;
N_248 <= CPI_M_PC_INTERNAL_15;
N_249 <= CPI_M_PC_INTERNAL_16;
N_250 <= CPI_M_PC_INTERNAL_17;
N_251 <= CPI_M_PC_INTERNAL_18;
N_252 <= CPI_M_PC_INTERNAL_19;
N_253 <= CPI_M_PC_INTERNAL_20;
N_254 <= CPI_M_PC_INTERNAL_21;
N_255 <= CPI_M_PC_INTERNAL_22;
N_256 <= CPI_M_PC_INTERNAL_23;
N_257 <= CPI_M_PC_INTERNAL_24;
N_258 <= CPI_M_PC_INTERNAL_25;
N_259 <= CPI_M_PC_INTERNAL_26;
N_260 <= CPI_M_PC_INTERNAL_27;
N_261 <= CPI_M_PC_INTERNAL_28;
N_262 <= CPI_M_PC_INTERNAL_29;
N_263 <= CPI_M_PC_INTERNAL_30;
N_264 <= CPI_M_INST_INTERNAL;
N_265 <= CPI_M_INST_INTERNAL_0;
N_266 <= CPI_M_INST_INTERNAL_1;
N_267 <= CPI_M_INST_INTERNAL_2;
N_268 <= CPI_M_INST_INTERNAL_3;
N_269 <= CPI_M_INST_INTERNAL_4;
N_270 <= CPI_M_INST_INTERNAL_5;
N_271 <= CPI_M_INST_INTERNAL_6;
N_272 <= CPI_M_INST_INTERNAL_7;
N_273 <= CPI_M_INST_INTERNAL_8;
N_274 <= CPI_M_INST_INTERNAL_9;
N_275 <= CPI_M_INST_INTERNAL_10;
N_276 <= CPI_M_INST_INTERNAL_11;
N_277 <= CPI_M_INST_INTERNAL_12;
N_278 <= CPI_M_INST_INTERNAL_13;
N_279 <= CPI_M_INST_INTERNAL_14;
N_280 <= CPI_M_INST_INTERNAL_15;
N_281 <= CPI_M_INST_INTERNAL_16;
N_282 <= CPI_M_INST_INTERNAL_17;
N_283 <= CPI_M_INST_INTERNAL_18;
N_284 <= CPI_M_INST_INTERNAL_19;
N_285 <= CPI_M_INST_INTERNAL_20;
N_286 <= CPI_M_INST_INTERNAL_21;
N_287 <= CPI_M_INST_INTERNAL_22;
N_288 <= CPI_M_INST_INTERNAL_23;
N_289 <= CPI_M_INST_INTERNAL_24;
N_290 <= CPI_M_INST_INTERNAL_25;
N_291 <= CPI_M_INST_INTERNAL_26;
N_292 <= CPI_M_INST_INTERNAL_27;
N_293 <= CPI_M_INST_INTERNAL_28;
N_294 <= CPI_M_INST_INTERNAL_29;
N_295 <= CPI_M_INST_INTERNAL_30;
N_296 <= CPI_M_CNT_INTERNAL;
N_297 <= CPI_M_CNT_INTERNAL_0;
N_298 <= CPI_M_TRAP_INTERNAL;
N_299 <= CPI_M_ANNUL_INTERNAL;
N_300 <= CPI_M_PV_INTERNAL;
N_301 <= CPI_X_PC_INTERNAL;
N_302 <= CPI_X_PC_INTERNAL_0;
N_303 <= CPI_X_PC_INTERNAL_1;
N_304 <= CPI_X_PC_INTERNAL_2;
N_305 <= CPI_X_PC_INTERNAL_3;
N_306 <= CPI_X_PC_INTERNAL_4;
N_307 <= CPI_X_PC_INTERNAL_5;
N_308 <= CPI_X_PC_INTERNAL_6;
N_309 <= CPI_X_PC_INTERNAL_7;
N_310 <= CPI_X_PC_INTERNAL_8;
N_311 <= CPI_X_PC_INTERNAL_9;
N_312 <= CPI_X_PC_INTERNAL_10;
N_313 <= CPI_X_PC_INTERNAL_11;
N_314 <= CPI_X_PC_INTERNAL_12;
N_315 <= CPI_X_PC_INTERNAL_13;
N_316 <= CPI_X_PC_INTERNAL_14;
N_317 <= CPI_X_PC_INTERNAL_15;
N_318 <= CPI_X_PC_INTERNAL_16;
N_319 <= CPI_X_PC_INTERNAL_17;
N_320 <= CPI_X_PC_INTERNAL_18;
N_321 <= CPI_X_PC_INTERNAL_19;
N_322 <= CPI_X_PC_INTERNAL_20;
N_323 <= CPI_X_PC_INTERNAL_21;
N_324 <= CPI_X_PC_INTERNAL_22;
N_325 <= CPI_X_PC_INTERNAL_23;
N_326 <= CPI_X_PC_INTERNAL_24;
N_327 <= CPI_X_PC_INTERNAL_25;
N_328 <= CPI_X_PC_INTERNAL_26;
N_329 <= CPI_X_PC_INTERNAL_27;
N_330 <= CPI_X_PC_INTERNAL_28;
N_331 <= CPI_X_PC_INTERNAL_29;
N_332 <= CPI_X_PC_INTERNAL_30;
N_333 <= CPI_X_INST_INTERNAL;
N_334 <= CPI_X_INST_INTERNAL_0;
N_335 <= CPI_X_INST_INTERNAL_1;
N_336 <= CPI_X_INST_INTERNAL_2;
N_337 <= CPI_X_INST_INTERNAL_3;
N_338 <= CPI_X_INST_INTERNAL_4;
N_339 <= CPI_X_INST_INTERNAL_5;
N_340 <= CPI_X_INST_INTERNAL_6;
N_341 <= CPI_X_INST_INTERNAL_7;
N_342 <= CPI_X_INST_INTERNAL_8;
N_343 <= CPI_X_INST_INTERNAL_9;
N_344 <= CPI_X_INST_INTERNAL_10;
N_345 <= CPI_X_INST_INTERNAL_11;
N_346 <= CPI_X_INST_INTERNAL_12;
N_347 <= CPI_X_INST_INTERNAL_13;
N_348 <= CPI_X_INST_INTERNAL_14;
N_349 <= CPI_X_INST_INTERNAL_15;
N_350 <= CPI_X_INST_INTERNAL_16;
N_351 <= CPI_X_INST_INTERNAL_17;
N_352 <= CPI_X_INST_INTERNAL_18;
N_353 <= CPI_X_INST_INTERNAL_19;
N_354 <= CPI_X_INST_INTERNAL_20;
N_355 <= CPI_X_INST_INTERNAL_21;
N_356 <= CPI_X_INST_INTERNAL_22;
N_357 <= CPI_X_INST_INTERNAL_23;
N_358 <= CPI_X_INST_INTERNAL_24;
N_359 <= CPI_X_INST_INTERNAL_25;
N_360 <= CPI_X_INST_INTERNAL_26;
N_361 <= CPI_X_INST_INTERNAL_27;
N_362 <= CPI_X_INST_INTERNAL_28;
N_363 <= CPI_X_INST_INTERNAL_29;
N_364 <= CPI_X_INST_INTERNAL_30;
N_365 <= CPI_X_CNT_INTERNAL;
N_366 <= CPI_X_CNT_INTERNAL_0;
N_367 <= CPI_X_TRAP_INTERNAL;
N_368 <= CPI_X_ANNUL_INTERNAL;
N_369 <= CPI_X_PV_INTERNAL;
N_370 <= CPI_LDDATA_INTERNAL;
N_371 <= CPI_LDDATA_INTERNAL_0;
N_372 <= CPI_LDDATA_INTERNAL_1;
N_373 <= CPI_LDDATA_INTERNAL_2;
N_374 <= CPI_LDDATA_INTERNAL_3;
N_375 <= CPI_LDDATA_INTERNAL_4;
N_376 <= CPI_LDDATA_INTERNAL_5;
N_377 <= CPI_LDDATA_INTERNAL_6;
N_378 <= CPI_LDDATA_INTERNAL_7;
N_379 <= CPI_LDDATA_INTERNAL_8;
N_380 <= CPI_LDDATA_INTERNAL_9;
N_381 <= CPI_LDDATA_INTERNAL_10;
N_382 <= CPI_LDDATA_INTERNAL_11;
N_383 <= CPI_LDDATA_INTERNAL_12;
N_384 <= CPI_LDDATA_INTERNAL_13;
N_385 <= CPI_LDDATA_INTERNAL_14;
N_386 <= CPI_LDDATA_INTERNAL_15;
N_387 <= CPI_LDDATA_INTERNAL_16;
N_388 <= CPI_LDDATA_INTERNAL_17;
N_389 <= CPI_LDDATA_INTERNAL_18;
N_390 <= CPI_LDDATA_INTERNAL_19;
N_391 <= CPI_LDDATA_INTERNAL_20;
N_392 <= CPI_LDDATA_INTERNAL_21;
N_393 <= CPI_LDDATA_INTERNAL_22;
N_394 <= CPI_LDDATA_INTERNAL_23;
N_395 <= CPI_LDDATA_INTERNAL_24;
N_396 <= CPI_LDDATA_INTERNAL_25;
N_397 <= CPI_LDDATA_INTERNAL_26;
N_398 <= CPI_LDDATA_INTERNAL_27;
N_399 <= CPI_LDDATA_INTERNAL_28;
N_400 <= CPI_LDDATA_INTERNAL_29;
N_401 <= CPI_LDDATA_INTERNAL_30;
N_402 <= CPI_DBG_ENABLE_INTERNAL;
N_403 <= CPI_DBG_WRITE_INTERNAL;
N_404 <= CPI_DBG_FSR_INTERNAL;
N_405 <= CPI_DBG_ADDR_INTERNAL;
N_406 <= CPI_DBG_ADDR_INTERNAL_0;
N_407 <= CPI_DBG_ADDR_INTERNAL_1;
N_408 <= CPI_DBG_ADDR_INTERNAL_2;
N_409 <= CPI_DBG_ADDR_INTERNAL_3;
N_410 <= CPI_DBG_DATA_INTERNAL;
N_411 <= CPI_DBG_DATA_INTERNAL_0;
N_412 <= CPI_DBG_DATA_INTERNAL_1;
N_413 <= CPI_DBG_DATA_INTERNAL_2;
N_414 <= CPI_DBG_DATA_INTERNAL_3;
N_415 <= CPI_DBG_DATA_INTERNAL_4;
N_416 <= CPI_DBG_DATA_INTERNAL_5;
N_417 <= CPI_DBG_DATA_INTERNAL_6;
N_418 <= CPI_DBG_DATA_INTERNAL_7;
N_419 <= CPI_DBG_DATA_INTERNAL_8;
N_420 <= CPI_DBG_DATA_INTERNAL_9;
N_421 <= CPI_DBG_DATA_INTERNAL_10;
N_422 <= CPI_DBG_DATA_INTERNAL_11;
N_423 <= CPI_DBG_DATA_INTERNAL_12;
N_424 <= CPI_DBG_DATA_INTERNAL_13;
N_425 <= CPI_DBG_DATA_INTERNAL_14;
N_426 <= CPI_DBG_DATA_INTERNAL_15;
N_427 <= CPI_DBG_DATA_INTERNAL_16;
N_428 <= CPI_DBG_DATA_INTERNAL_17;
N_429 <= CPI_DBG_DATA_INTERNAL_18;
N_430 <= CPI_DBG_DATA_INTERNAL_19;
N_431 <= CPI_DBG_DATA_INTERNAL_20;
N_432 <= CPI_DBG_DATA_INTERNAL_21;
N_433 <= CPI_DBG_DATA_INTERNAL_22;
N_434 <= CPI_DBG_DATA_INTERNAL_23;
N_435 <= CPI_DBG_DATA_INTERNAL_24;
N_436 <= CPI_DBG_DATA_INTERNAL_25;
N_437 <= CPI_DBG_DATA_INTERNAL_26;
N_438 <= CPI_DBG_DATA_INTERNAL_27;
N_439 <= CPI_DBG_DATA_INTERNAL_28;
N_440 <= CPI_DBG_DATA_INTERNAL_29;
N_441 <= CPI_DBG_DATA_INTERNAL_30;
N_0 <= CPO_DATAZ(0);
N_1_72 <= CPO_DATAZ(1);
N_2_0 <= CPO_DATAZ(2);
N_3_0 <= CPO_DATAZ(3);
N_4_0 <= CPO_DATAZ(4);
N_5_0 <= CPO_DATAZ(5);
N_6_0 <= CPO_DATAZ(6);
N_7_0 <= CPO_DATAZ(7);
N_8_0 <= CPO_DATAZ(8);
N_9_0 <= CPO_DATAZ(9);
N_10_1 <= CPO_DATAZ(10);
N_11_2 <= CPO_DATAZ(11);
N_12_1 <= CPO_DATAZ(12);
N_13_1 <= CPO_DATAZ(13);
N_14_0 <= CPO_DATAZ(14);
N_15_0 <= CPO_DATAZ(15);
N_16_0 <= CPO_DATAZ(16);
N_17_0 <= CPO_DATAZ(17);
N_18_0 <= CPO_DATAZ(18);
N_19_0 <= CPO_DATAZ(19);
N_20_0 <= CPO_DATAZ(20);
N_21_0 <= CPO_DATAZ(21);
N_22_0 <= CPO_DATAZ(22);
N_23_0 <= CPO_DATAZ(23);
N_24_0 <= CPO_DATAZ(24);
N_25_0 <= CPO_DATAZ(25);
N_26_0 <= CPO_DATAZ(26);
N_27_0 <= CPO_DATAZ(27);
N_28_0 <= CPO_DATAZ(28);
N_29_0 <= CPO_DATAZ(29);
N_30_0 <= CPO_DATAZ(30);
N_31_0 <= CPO_DATAZ(31);
N_32_0 <= CPO_EXCZ;
N_33_0 <= CPO_CCZ(0);
N_34_0 <= CPO_CCZ(1);
N_35_0 <= CPO_CCVZ;
N_36_0 <= CPO_LDLOCKZ;
N_37_0 <= CPO_HOLDNZ;
N_38_0 <= CPO_DBG_DATAZ(0);
N_39_0 <= CPO_DBG_DATAZ(1);
N_40_0 <= CPO_DBG_DATAZ(2);
N_41_0 <= CPO_DBG_DATAZ(3);
N_42_0 <= CPO_DBG_DATAZ(4);
N_43_0 <= CPO_DBG_DATAZ(5);
N_44_0 <= CPO_DBG_DATAZ(6);
N_45_0 <= CPO_DBG_DATAZ(7);
N_46_0 <= CPO_DBG_DATAZ(8);
N_47_0 <= CPO_DBG_DATAZ(9);
N_48_0 <= CPO_DBG_DATAZ(10);
N_49_0 <= CPO_DBG_DATAZ(11);
N_50_0 <= CPO_DBG_DATAZ(12);
N_51_0 <= CPO_DBG_DATAZ(13);
N_52_0 <= CPO_DBG_DATAZ(14);
N_53_0 <= CPO_DBG_DATAZ(15);
N_54_0 <= CPO_DBG_DATAZ(16);
N_55_0 <= CPO_DBG_DATAZ(17);
N_56_0 <= CPO_DBG_DATAZ(18);
N_57_0 <= CPO_DBG_DATAZ(19);
N_58_0 <= CPO_DBG_DATAZ(20);
N_59_0 <= CPO_DBG_DATAZ(21);
N_60_0 <= CPO_DBG_DATAZ(22);
N_61_0 <= CPO_DBG_DATAZ(23);
N_62_0 <= CPO_DBG_DATAZ(24);
N_63_0 <= CPO_DBG_DATAZ(25);
N_64_0 <= CPO_DBG_DATAZ(26);
N_65_0 <= CPO_DBG_DATAZ(27);
N_66_0 <= CPO_DBG_DATAZ(28);
N_67_0 <= CPO_DBG_DATAZ(29);
N_68_0 <= CPO_DBG_DATAZ(30);
N_69_0 <= CPO_DBG_DATAZ(31);
N_70_0 <= RFI2_RD1ADDRZ(0);
N_71_0 <= RFI2_RD1ADDRZ(1);
N_72_0 <= RFI2_RD1ADDRZ(2);
N_73_0 <= RFI2_RD1ADDRZ(3);
N_74_0 <= RFI2_RD2ADDRZ(0);
N_75_0 <= RFI2_RD2ADDRZ(1);
N_76_0 <= RFI2_RD2ADDRZ(2);
N_77_0 <= RFI2_RD2ADDRZ(3);
N_78_0 <= RFI2_WRADDRZ(0);
N_79_0 <= RFI2_WRADDRZ(1);
N_80_0 <= RFI2_WRADDRZ(2);
N_81_0 <= RFI2_WRADDRZ(3);
N_82_0 <= RFI1_WRDATAZ(0);
N_83_0 <= RFI1_WRDATAZ(1);
N_84_0 <= RFI1_WRDATAZ(2);
N_85_0 <= RFI1_WRDATAZ(3);
N_86_0 <= RFI1_WRDATAZ(4);
N_87_0 <= RFI1_WRDATAZ(5);
N_88_0 <= RFI1_WRDATAZ(6);
N_89_0 <= RFI1_WRDATAZ(7);
N_90_0 <= RFI1_WRDATAZ(8);
N_91_0 <= RFI1_WRDATAZ(9);
N_92_0 <= RFI1_WRDATAZ(10);
N_93_0 <= RFI1_WRDATAZ(11);
N_94_0 <= RFI1_WRDATAZ(12);
N_95_0 <= RFI1_WRDATAZ(13);
N_96_0 <= RFI1_WRDATAZ(14);
N_97_0 <= RFI1_WRDATAZ(15);
N_98_0 <= RFI1_WRDATAZ(16);
N_99_0 <= RFI1_WRDATAZ(17);
N_100_0 <= RFI1_WRDATAZ(18);
N_101_0 <= RFI1_WRDATAZ(19);
N_102_0 <= RFI1_WRDATAZ(20);
N_103_0 <= RFI1_WRDATAZ(21);
N_104_0 <= RFI1_WRDATAZ(22);
N_105_0 <= RFI1_WRDATAZ(23);
N_106_0 <= RFI1_WRDATAZ(24);
N_107_0 <= RFI1_WRDATAZ(25);
N_108_0 <= RFI1_WRDATAZ(26);
N_109_0 <= RFI1_WRDATAZ(27);
N_110_0 <= RFI1_WRDATAZ(28);
N_111_0 <= RFI1_WRDATAZ(29);
N_112_0 <= RFI1_WRDATAZ(30);
N_113_0 <= RFI1_WRDATAZ(31);
N_114_0 <= RFI1_REN1Z;
N_115_0 <= RFI1_REN2Z;
N_116_0 <= RFI1_WRENZ;
N_117_0 <= RFI2_RD1ADDRZ(0);
N_118_0 <= RFI2_RD1ADDRZ(1);
N_119_0 <= RFI2_RD1ADDRZ(2);
N_120_0 <= RFI2_RD1ADDRZ(3);
N_121_0 <= RFI2_RD2ADDRZ(0);
N_122_0 <= RFI2_RD2ADDRZ(1);
N_123_0 <= RFI2_RD2ADDRZ(2);
N_124_0 <= RFI2_RD2ADDRZ(3);
N_125_0 <= RFI2_WRADDRZ(0);
N_126_0 <= RFI2_WRADDRZ(1);
N_127_0 <= RFI2_WRADDRZ(2);
N_128_0 <= RFI2_WRADDRZ(3);
N_129_0 <= RFI2_WRDATAZ(0);
N_130_0 <= RFI2_WRDATAZ(1);
N_131_0 <= RFI2_WRDATAZ(2);
N_132_0 <= RFI2_WRDATAZ(3);
N_133_0 <= RFI2_WRDATAZ(4);
N_134_0 <= RFI2_WRDATAZ(5);
N_135_0 <= RFI2_WRDATAZ(6);
N_136_0 <= RFI2_WRDATAZ(7);
N_137_0 <= RFI2_WRDATAZ(8);
N_138_0 <= RFI2_WRDATAZ(9);
N_139_0 <= RFI2_WRDATAZ(10);
N_140_0 <= RFI2_WRDATAZ(11);
N_141_0 <= RFI2_WRDATAZ(12);
N_142_0 <= RFI2_WRDATAZ(13);
N_143_0 <= RFI2_WRDATAZ(14);
N_144_0 <= RFI2_WRDATAZ(15);
N_145_0 <= RFI2_WRDATAZ(16);
N_146_0 <= RFI2_WRDATAZ(17);
N_147_0 <= RFI2_WRDATAZ(18);
N_148_0 <= RFI2_WRDATAZ(19);
N_149_0 <= RFI2_WRDATAZ(20);
N_150_0 <= RFI2_WRDATAZ(21);
N_151_0 <= RFI2_WRDATAZ(22);
N_152_0 <= RFI2_WRDATAZ(23);
N_153_0 <= RFI2_WRDATAZ(24);
N_154_0 <= RFI2_WRDATAZ(25);
N_155_0 <= RFI2_WRDATAZ(26);
N_156_0 <= RFI2_WRDATAZ(27);
N_157_0 <= RFI2_WRDATAZ(28);
N_158_0 <= RFI2_WRDATAZ(29);
N_159_0 <= RFI2_WRDATAZ(30);
N_160_0 <= RFI2_WRDATAZ(31);
N_161_0 <= RFI2_REN1Z;
N_162_0 <= RFI2_REN2Z;
N_163_0 <= RFI2_WRENZ;
N_606 <= RFO1_DATA1_INTERNAL;
N_607 <= RFO1_DATA1_INTERNAL_0;
N_608 <= RFO1_DATA1_INTERNAL_1;
N_609 <= RFO1_DATA1_INTERNAL_2;
N_610 <= RFO1_DATA1_INTERNAL_3;
N_611 <= RFO1_DATA1_INTERNAL_4;
N_612 <= RFO1_DATA1_INTERNAL_5;
N_613 <= RFO1_DATA1_INTERNAL_6;
N_614 <= RFO1_DATA1_INTERNAL_7;
N_615 <= RFO1_DATA1_INTERNAL_8;
N_616 <= RFO1_DATA1_INTERNAL_9;
N_617 <= RFO1_DATA1_INTERNAL_10;
N_618 <= RFO1_DATA1_INTERNAL_11;
N_619 <= RFO1_DATA1_INTERNAL_12;
N_620 <= RFO1_DATA1_INTERNAL_13;
N_621 <= RFO1_DATA1_INTERNAL_14;
N_622 <= RFO1_DATA1_INTERNAL_15;
N_623 <= RFO1_DATA1_INTERNAL_16;
N_624 <= RFO1_DATA1_INTERNAL_17;
N_625 <= RFO1_DATA1_INTERNAL_18;
N_626 <= RFO1_DATA1_INTERNAL_19;
N_627 <= RFO1_DATA1_INTERNAL_20;
N_628 <= RFO1_DATA1_INTERNAL_21;
N_629 <= RFO1_DATA1_INTERNAL_22;
N_630 <= RFO1_DATA1_INTERNAL_23;
N_631 <= RFO1_DATA1_INTERNAL_24;
N_632 <= RFO1_DATA1_INTERNAL_25;
N_633 <= RFO1_DATA1_INTERNAL_26;
N_634 <= RFO1_DATA1_INTERNAL_27;
N_635 <= RFO1_DATA1_INTERNAL_28;
N_636 <= RFO1_DATA1_INTERNAL_29;
N_637 <= RFO1_DATA1_INTERNAL_30;
N_638 <= RFO1_DATA2_INTERNAL;
N_639 <= RFO1_DATA2_INTERNAL_0;
N_640 <= RFO1_DATA2_INTERNAL_1;
N_641 <= RFO1_DATA2_INTERNAL_2;
N_642 <= RFO1_DATA2_INTERNAL_3;
N_643 <= RFO1_DATA2_INTERNAL_4;
N_644 <= RFO1_DATA2_INTERNAL_5;
N_645 <= RFO1_DATA2_INTERNAL_6;
N_646 <= RFO1_DATA2_INTERNAL_7;
N_647 <= RFO1_DATA2_INTERNAL_8;
N_648 <= RFO1_DATA2_INTERNAL_9;
N_649 <= RFO1_DATA2_INTERNAL_10;
N_650 <= RFO1_DATA2_INTERNAL_11;
N_651 <= RFO1_DATA2_INTERNAL_12;
N_652 <= RFO1_DATA2_INTERNAL_13;
N_653 <= RFO1_DATA2_INTERNAL_14;
N_654 <= RFO1_DATA2_INTERNAL_15;
N_655 <= RFO1_DATA2_INTERNAL_16;
N_656 <= RFO1_DATA2_INTERNAL_17;
N_657 <= RFO1_DATA2_INTERNAL_18;
N_658 <= RFO1_DATA2_INTERNAL_19;
N_659 <= RFO1_DATA2_INTERNAL_20;
N_660 <= RFO1_DATA2_INTERNAL_21;
N_661 <= RFO1_DATA2_INTERNAL_22;
N_662 <= RFO1_DATA2_INTERNAL_23;
N_663 <= RFO1_DATA2_INTERNAL_24;
N_664 <= RFO1_DATA2_INTERNAL_25;
N_665 <= RFO1_DATA2_INTERNAL_26;
N_666 <= RFO1_DATA2_INTERNAL_27;
N_667 <= RFO1_DATA2_INTERNAL_28;
N_668 <= RFO1_DATA2_INTERNAL_29;
N_669 <= RFO1_DATA2_INTERNAL_30;
N_670 <= RFO2_DATA1_INTERNAL;
N_671 <= RFO2_DATA1_INTERNAL_0;
N_672 <= RFO2_DATA1_INTERNAL_1;
N_673 <= RFO2_DATA1_INTERNAL_2;
N_674 <= RFO2_DATA1_INTERNAL_3;
N_675 <= RFO2_DATA1_INTERNAL_4;
N_676 <= RFO2_DATA1_INTERNAL_5;
N_677 <= RFO2_DATA1_INTERNAL_6;
N_678 <= RFO2_DATA1_INTERNAL_7;
N_679 <= RFO2_DATA1_INTERNAL_8;
N_680 <= RFO2_DATA1_INTERNAL_9;
N_681 <= RFO2_DATA1_INTERNAL_10;
N_682 <= RFO2_DATA1_INTERNAL_11;
N_683 <= RFO2_DATA1_INTERNAL_12;
N_684 <= RFO2_DATA1_INTERNAL_13;
N_685 <= RFO2_DATA1_INTERNAL_14;
N_686 <= RFO2_DATA1_INTERNAL_15;
N_687 <= RFO2_DATA1_INTERNAL_16;
N_688 <= RFO2_DATA1_INTERNAL_17;
N_689 <= RFO2_DATA1_INTERNAL_18;
N_690 <= RFO2_DATA1_INTERNAL_19;
N_691 <= RFO2_DATA1_INTERNAL_20;
N_692 <= RFO2_DATA1_INTERNAL_21;
N_693 <= RFO2_DATA1_INTERNAL_22;
N_694 <= RFO2_DATA1_INTERNAL_23;
N_695 <= RFO2_DATA1_INTERNAL_24;
N_696 <= RFO2_DATA1_INTERNAL_25;
N_697 <= RFO2_DATA1_INTERNAL_26;
N_698 <= RFO2_DATA1_INTERNAL_27;
N_699 <= RFO2_DATA1_INTERNAL_28;
N_700 <= RFO2_DATA1_INTERNAL_29;
N_701 <= RFO2_DATA1_INTERNAL_30;
N_702 <= RFO2_DATA2_INTERNAL;
N_703 <= RFO2_DATA2_INTERNAL_0;
N_704 <= RFO2_DATA2_INTERNAL_1;
N_705 <= RFO2_DATA2_INTERNAL_2;
N_706 <= RFO2_DATA2_INTERNAL_3;
N_707 <= RFO2_DATA2_INTERNAL_4;
N_708 <= RFO2_DATA2_INTERNAL_5;
N_709 <= RFO2_DATA2_INTERNAL_6;
N_710 <= RFO2_DATA2_INTERNAL_7;
N_711 <= RFO2_DATA2_INTERNAL_8;
N_712 <= RFO2_DATA2_INTERNAL_9;
N_713 <= RFO2_DATA2_INTERNAL_10;
N_714 <= RFO2_DATA2_INTERNAL_11;
N_715 <= RFO2_DATA2_INTERNAL_12;
N_716 <= RFO2_DATA2_INTERNAL_13;
N_717 <= RFO2_DATA2_INTERNAL_14;
N_718 <= RFO2_DATA2_INTERNAL_15;
N_719 <= RFO2_DATA2_INTERNAL_16;
N_720 <= RFO2_DATA2_INTERNAL_17;
N_721 <= RFO2_DATA2_INTERNAL_18;
N_722 <= RFO2_DATA2_INTERNAL_19;
N_723 <= RFO2_DATA2_INTERNAL_20;
N_724 <= RFO2_DATA2_INTERNAL_21;
N_725 <= RFO2_DATA2_INTERNAL_22;
N_726 <= RFO2_DATA2_INTERNAL_23;
N_727 <= RFO2_DATA2_INTERNAL_24;
N_728 <= RFO2_DATA2_INTERNAL_25;
N_729 <= RFO2_DATA2_INTERNAL_26;
N_730 <= RFO2_DATA2_INTERNAL_27;
N_731 <= RFO2_DATA2_INTERNAL_28;
N_732 <= RFO2_DATA2_INTERNAL_29;
N_733 <= RFO2_DATA2_INTERNAL_30;
\GRLFPC2_0.COMB.V.A.AFQ_1_I\ <= not \GRLFPC2_0.COMB.V.A.AFQ_1\;
\GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4_I\ <= not \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_1_SN_M4\;
\GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3_I\ <= not \GRLFPC2_0.GRFPUL_GEN0.GRFPULITE0.RIN.DPATH_SN_M3\;
\GRLFPC2_0.COMB.UN2_HOLDN_0_A2_I\ <= not \GRLFPC2_0.COMB.UN2_HOLDN_0_A2\;
\GRLFPC2_0.FPI.LDOP_I\ <= not \GRLFPC2_0.FPI.LDOP\;
cpo_data(0) <= N_0;
cpo_data(1) <= N_1_72;
cpo_data(2) <= N_2_0;
cpo_data(3) <= N_3_0;
cpo_data(4) <= N_4_0;
cpo_data(5) <= N_5_0;
cpo_data(6) <= N_6_0;
cpo_data(7) <= N_7_0;
cpo_data(8) <= N_8_0;
cpo_data(9) <= N_9_0;
cpo_data(10) <= N_10_1;
cpo_data(11) <= N_11_2;
cpo_data(12) <= N_12_1;
cpo_data(13) <= N_13_1;
cpo_data(14) <= N_14_0;
cpo_data(15) <= N_15_0;
cpo_data(16) <= N_16_0;
cpo_data(17) <= N_17_0;
cpo_data(18) <= N_18_0;
cpo_data(19) <= N_19_0;
cpo_data(20) <= N_20_0;
cpo_data(21) <= N_21_0;
cpo_data(22) <= N_22_0;
cpo_data(23) <= N_23_0;
cpo_data(24) <= N_24_0;
cpo_data(25) <= N_25_0;
cpo_data(26) <= N_26_0;
cpo_data(27) <= N_27_0;
cpo_data(28) <= N_28_0;
cpo_data(29) <= N_29_0;
cpo_data(30) <= N_30_0;
cpo_data(31) <= N_31_0;
cpo_exc <= N_32_0;
cpo_cc(0) <= N_33_0;
cpo_cc(1) <= N_34_0;
cpo_ccv <= N_35_0;
cpo_ldlock <= N_36_0;
cpo_holdn <= N_37_0;
cpo_dbg_data(0) <= N_38_0;
cpo_dbg_data(1) <= N_39_0;
cpo_dbg_data(2) <= N_40_0;
cpo_dbg_data(3) <= N_41_0;
cpo_dbg_data(4) <= N_42_0;
cpo_dbg_data(5) <= N_43_0;
cpo_dbg_data(6) <= N_44_0;
cpo_dbg_data(7) <= N_45_0;
cpo_dbg_data(8) <= N_46_0;
cpo_dbg_data(9) <= N_47_0;
cpo_dbg_data(10) <= N_48_0;
cpo_dbg_data(11) <= N_49_0;
cpo_dbg_data(12) <= N_50_0;
cpo_dbg_data(13) <= N_51_0;
cpo_dbg_data(14) <= N_52_0;
cpo_dbg_data(15) <= N_53_0;
cpo_dbg_data(16) <= N_54_0;
cpo_dbg_data(17) <= N_55_0;
cpo_dbg_data(18) <= N_56_0;
cpo_dbg_data(19) <= N_57_0;
cpo_dbg_data(20) <= N_58_0;
cpo_dbg_data(21) <= N_59_0;
cpo_dbg_data(22) <= N_60_0;
cpo_dbg_data(23) <= N_61_0;
cpo_dbg_data(24) <= N_62_0;
cpo_dbg_data(25) <= N_63_0;
cpo_dbg_data(26) <= N_64_0;
cpo_dbg_data(27) <= N_65_0;
cpo_dbg_data(28) <= N_66_0;
cpo_dbg_data(29) <= N_67_0;
cpo_dbg_data(30) <= N_68_0;
cpo_dbg_data(31) <= N_69_0;
rfi1_rd1addr(0) <= N_70_0;
rfi1_rd1addr(1) <= N_71_0;
rfi1_rd1addr(2) <= N_72_0;
rfi1_rd1addr(3) <= N_73_0;
rfi1_rd2addr(0) <= N_74_0;
rfi1_rd2addr(1) <= N_75_0;
rfi1_rd2addr(2) <= N_76_0;
rfi1_rd2addr(3) <= N_77_0;
rfi1_wraddr(0) <= N_78_0;
rfi1_wraddr(1) <= N_79_0;
rfi1_wraddr(2) <= N_80_0;
rfi1_wraddr(3) <= N_81_0;
rfi1_wrdata(0) <= N_82_0;
rfi1_wrdata(1) <= N_83_0;
rfi1_wrdata(2) <= N_84_0;
rfi1_wrdata(3) <= N_85_0;
rfi1_wrdata(4) <= N_86_0;
rfi1_wrdata(5) <= N_87_0;
rfi1_wrdata(6) <= N_88_0;
rfi1_wrdata(7) <= N_89_0;
rfi1_wrdata(8) <= N_90_0;
rfi1_wrdata(9) <= N_91_0;
rfi1_wrdata(10) <= N_92_0;
rfi1_wrdata(11) <= N_93_0;
rfi1_wrdata(12) <= N_94_0;
rfi1_wrdata(13) <= N_95_0;
rfi1_wrdata(14) <= N_96_0;
rfi1_wrdata(15) <= N_97_0;
rfi1_wrdata(16) <= N_98_0;
rfi1_wrdata(17) <= N_99_0;
rfi1_wrdata(18) <= N_100_0;
rfi1_wrdata(19) <= N_101_0;
rfi1_wrdata(20) <= N_102_0;
rfi1_wrdata(21) <= N_103_0;
rfi1_wrdata(22) <= N_104_0;
rfi1_wrdata(23) <= N_105_0;
rfi1_wrdata(24) <= N_106_0;
rfi1_wrdata(25) <= N_107_0;
rfi1_wrdata(26) <= N_108_0;
rfi1_wrdata(27) <= N_109_0;
rfi1_wrdata(28) <= N_110_0;
rfi1_wrdata(29) <= N_111_0;
rfi1_wrdata(30) <= N_112_0;
rfi1_wrdata(31) <= N_113_0;
rfi1_ren1 <= N_114_0;
rfi1_ren2 <= N_115_0;
rfi1_wren <= N_116_0;
rfi2_rd1addr(0) <= N_117_0;
rfi2_rd1addr(1) <= N_118_0;
rfi2_rd1addr(2) <= N_119_0;
rfi2_rd1addr(3) <= N_120_0;
rfi2_rd2addr(0) <= N_121_0;
rfi2_rd2addr(1) <= N_122_0;
rfi2_rd2addr(2) <= N_123_0;
rfi2_rd2addr(3) <= N_124_0;
rfi2_wraddr(0) <= N_125_0;
rfi2_wraddr(1) <= N_126_0;
rfi2_wraddr(2) <= N_127_0;
rfi2_wraddr(3) <= N_128_0;
rfi2_wrdata(0) <= N_129_0;
rfi2_wrdata(1) <= N_130_0;
rfi2_wrdata(2) <= N_131_0;
rfi2_wrdata(3) <= N_132_0;
rfi2_wrdata(4) <= N_133_0;
rfi2_wrdata(5) <= N_134_0;
rfi2_wrdata(6) <= N_135_0;
rfi2_wrdata(7) <= N_136_0;
rfi2_wrdata(8) <= N_137_0;
rfi2_wrdata(9) <= N_138_0;
rfi2_wrdata(10) <= N_139_0;
rfi2_wrdata(11) <= N_140_0;
rfi2_wrdata(12) <= N_141_0;
rfi2_wrdata(13) <= N_142_0;
rfi2_wrdata(14) <= N_143_0;
rfi2_wrdata(15) <= N_144_0;
rfi2_wrdata(16) <= N_145_0;
rfi2_wrdata(17) <= N_146_0;
rfi2_wrdata(18) <= N_147_0;
rfi2_wrdata(19) <= N_148_0;
rfi2_wrdata(20) <= N_149_0;
rfi2_wrdata(21) <= N_150_0;
rfi2_wrdata(22) <= N_151_0;
rfi2_wrdata(23) <= N_152_0;
rfi2_wrdata(24) <= N_153_0;
rfi2_wrdata(25) <= N_154_0;
rfi2_wrdata(26) <= N_155_0;
rfi2_wrdata(27) <= N_156_0;
rfi2_wrdata(28) <= N_157_0;
rfi2_wrdata(29) <= N_158_0;
rfi2_wrdata(30) <= N_159_0;
rfi2_wrdata(31) <= N_160_0;
rfi2_ren1 <= N_161_0;
rfi2_ren2 <= N_162_0;
rfi2_wren <= N_163_0;
RST_INTERNAL <= rst;
CLK_INTERNAL <= clk;
HOLDN_INTERNAL <= holdn;
CPI_FLUSH_INTERNAL <= cpi_flush;
CPI_EXACK_INTERNAL <= cpi_exack;
CPI_A_RS1_INTERNAL <= cpi_a_rs1(0);
CPI_A_RS1_INTERNAL_0 <= cpi_a_rs1(1);
CPI_A_RS1_INTERNAL_1 <= cpi_a_rs1(2);
CPI_A_RS1_INTERNAL_2 <= cpi_a_rs1(3);
CPI_A_RS1_INTERNAL_3 <= cpi_a_rs1(4);
CPI_D_PC_INTERNAL <= cpi_d_pc(0);
CPI_D_PC_INTERNAL_0 <= cpi_d_pc(1);
CPI_D_PC_INTERNAL_1 <= cpi_d_pc(2);
CPI_D_PC_INTERNAL_2 <= cpi_d_pc(3);
CPI_D_PC_INTERNAL_3 <= cpi_d_pc(4);
CPI_D_PC_INTERNAL_4 <= cpi_d_pc(5);
CPI_D_PC_INTERNAL_5 <= cpi_d_pc(6);
CPI_D_PC_INTERNAL_6 <= cpi_d_pc(7);
CPI_D_PC_INTERNAL_7 <= cpi_d_pc(8);
CPI_D_PC_INTERNAL_8 <= cpi_d_pc(9);
CPI_D_PC_INTERNAL_9 <= cpi_d_pc(10);
CPI_D_PC_INTERNAL_10 <= cpi_d_pc(11);
CPI_D_PC_INTERNAL_11 <= cpi_d_pc(12);
CPI_D_PC_INTERNAL_12 <= cpi_d_pc(13);
CPI_D_PC_INTERNAL_13 <= cpi_d_pc(14);
CPI_D_PC_INTERNAL_14 <= cpi_d_pc(15);
CPI_D_PC_INTERNAL_15 <= cpi_d_pc(16);
CPI_D_PC_INTERNAL_16 <= cpi_d_pc(17);
CPI_D_PC_INTERNAL_17 <= cpi_d_pc(18);
CPI_D_PC_INTERNAL_18 <= cpi_d_pc(19);
CPI_D_PC_INTERNAL_19 <= cpi_d_pc(20);
CPI_D_PC_INTERNAL_20 <= cpi_d_pc(21);
CPI_D_PC_INTERNAL_21 <= cpi_d_pc(22);
CPI_D_PC_INTERNAL_22 <= cpi_d_pc(23);
CPI_D_PC_INTERNAL_23 <= cpi_d_pc(24);
CPI_D_PC_INTERNAL_24 <= cpi_d_pc(25);
CPI_D_PC_INTERNAL_25 <= cpi_d_pc(26);
CPI_D_PC_INTERNAL_26 <= cpi_d_pc(27);
CPI_D_PC_INTERNAL_27 <= cpi_d_pc(28);
CPI_D_PC_INTERNAL_28 <= cpi_d_pc(29);
CPI_D_PC_INTERNAL_29 <= cpi_d_pc(30);
CPI_D_PC_INTERNAL_30 <= cpi_d_pc(31);
CPI_D_INST_INTERNAL <= cpi_d_inst(0);
CPI_D_INST_INTERNAL_0 <= cpi_d_inst(1);
CPI_D_INST_INTERNAL_1 <= cpi_d_inst(2);
CPI_D_INST_INTERNAL_2 <= cpi_d_inst(3);
CPI_D_INST_INTERNAL_3 <= cpi_d_inst(4);
CPI_D_INST_INTERNAL_4 <= cpi_d_inst(5);
CPI_D_INST_INTERNAL_5 <= cpi_d_inst(6);
CPI_D_INST_INTERNAL_6 <= cpi_d_inst(7);
CPI_D_INST_INTERNAL_7 <= cpi_d_inst(8);
CPI_D_INST_INTERNAL_8 <= cpi_d_inst(9);
CPI_D_INST_INTERNAL_9 <= cpi_d_inst(10);
CPI_D_INST_INTERNAL_10 <= cpi_d_inst(11);
CPI_D_INST_INTERNAL_11 <= cpi_d_inst(12);
CPI_D_INST_INTERNAL_12 <= cpi_d_inst(13);
CPI_D_INST_INTERNAL_13 <= cpi_d_inst(14);
CPI_D_INST_INTERNAL_14 <= cpi_d_inst(15);
CPI_D_INST_INTERNAL_15 <= cpi_d_inst(16);
CPI_D_INST_INTERNAL_16 <= cpi_d_inst(17);
CPI_D_INST_INTERNAL_17 <= cpi_d_inst(18);
CPI_D_INST_INTERNAL_18 <= cpi_d_inst(19);
CPI_D_INST_INTERNAL_19 <= cpi_d_inst(20);
CPI_D_INST_INTERNAL_20 <= cpi_d_inst(21);
CPI_D_INST_INTERNAL_21 <= cpi_d_inst(22);
CPI_D_INST_INTERNAL_22 <= cpi_d_inst(23);
CPI_D_INST_INTERNAL_23 <= cpi_d_inst(24);
CPI_D_INST_INTERNAL_24 <= cpi_d_inst(25);
CPI_D_INST_INTERNAL_25 <= cpi_d_inst(26);
CPI_D_INST_INTERNAL_26 <= cpi_d_inst(27);
CPI_D_INST_INTERNAL_27 <= cpi_d_inst(28);
CPI_D_INST_INTERNAL_28 <= cpi_d_inst(29);
CPI_D_INST_INTERNAL_29 <= cpi_d_inst(30);
CPI_D_INST_INTERNAL_30 <= cpi_d_inst(31);
CPI_D_CNT_INTERNAL <= cpi_d_cnt(0);
CPI_D_CNT_INTERNAL_0 <= cpi_d_cnt(1);
CPI_D_TRAP_INTERNAL <= cpi_d_trap;
CPI_D_ANNUL_INTERNAL <= cpi_d_annul;
CPI_D_PV_INTERNAL <= cpi_d_pv;
CPI_A_PC_INTERNAL <= cpi_a_pc(0);
CPI_A_PC_INTERNAL_0 <= cpi_a_pc(1);
CPI_A_PC_INTERNAL_1 <= cpi_a_pc(2);
CPI_A_PC_INTERNAL_2 <= cpi_a_pc(3);
CPI_A_PC_INTERNAL_3 <= cpi_a_pc(4);
CPI_A_PC_INTERNAL_4 <= cpi_a_pc(5);
CPI_A_PC_INTERNAL_5 <= cpi_a_pc(6);
CPI_A_PC_INTERNAL_6 <= cpi_a_pc(7);
CPI_A_PC_INTERNAL_7 <= cpi_a_pc(8);
CPI_A_PC_INTERNAL_8 <= cpi_a_pc(9);
CPI_A_PC_INTERNAL_9 <= cpi_a_pc(10);
CPI_A_PC_INTERNAL_10 <= cpi_a_pc(11);
CPI_A_PC_INTERNAL_11 <= cpi_a_pc(12);
CPI_A_PC_INTERNAL_12 <= cpi_a_pc(13);
CPI_A_PC_INTERNAL_13 <= cpi_a_pc(14);
CPI_A_PC_INTERNAL_14 <= cpi_a_pc(15);
CPI_A_PC_INTERNAL_15 <= cpi_a_pc(16);
CPI_A_PC_INTERNAL_16 <= cpi_a_pc(17);
CPI_A_PC_INTERNAL_17 <= cpi_a_pc(18);
CPI_A_PC_INTERNAL_18 <= cpi_a_pc(19);
CPI_A_PC_INTERNAL_19 <= cpi_a_pc(20);
CPI_A_PC_INTERNAL_20 <= cpi_a_pc(21);
CPI_A_PC_INTERNAL_21 <= cpi_a_pc(22);
CPI_A_PC_INTERNAL_22 <= cpi_a_pc(23);
CPI_A_PC_INTERNAL_23 <= cpi_a_pc(24);
CPI_A_PC_INTERNAL_24 <= cpi_a_pc(25);
CPI_A_PC_INTERNAL_25 <= cpi_a_pc(26);
CPI_A_PC_INTERNAL_26 <= cpi_a_pc(27);
CPI_A_PC_INTERNAL_27 <= cpi_a_pc(28);
CPI_A_PC_INTERNAL_28 <= cpi_a_pc(29);
CPI_A_PC_INTERNAL_29 <= cpi_a_pc(30);
CPI_A_PC_INTERNAL_30 <= cpi_a_pc(31);
CPI_A_INST_INTERNAL <= cpi_a_inst(0);
CPI_A_INST_INTERNAL_0 <= cpi_a_inst(1);
CPI_A_INST_INTERNAL_1 <= cpi_a_inst(2);
CPI_A_INST_INTERNAL_2 <= cpi_a_inst(3);
CPI_A_INST_INTERNAL_3 <= cpi_a_inst(4);
CPI_A_INST_INTERNAL_4 <= cpi_a_inst(5);
CPI_A_INST_INTERNAL_5 <= cpi_a_inst(6);
CPI_A_INST_INTERNAL_6 <= cpi_a_inst(7);
CPI_A_INST_INTERNAL_7 <= cpi_a_inst(8);
CPI_A_INST_INTERNAL_8 <= cpi_a_inst(9);
CPI_A_INST_INTERNAL_9 <= cpi_a_inst(10);
CPI_A_INST_INTERNAL_10 <= cpi_a_inst(11);
CPI_A_INST_INTERNAL_11 <= cpi_a_inst(12);
CPI_A_INST_INTERNAL_12 <= cpi_a_inst(13);
CPI_A_INST_INTERNAL_13 <= cpi_a_inst(14);
CPI_A_INST_INTERNAL_14 <= cpi_a_inst(15);
CPI_A_INST_INTERNAL_15 <= cpi_a_inst(16);
CPI_A_INST_INTERNAL_16 <= cpi_a_inst(17);
CPI_A_INST_INTERNAL_17 <= cpi_a_inst(18);
CPI_A_INST_INTERNAL_18 <= cpi_a_inst(19);
CPI_A_INST_INTERNAL_19 <= cpi_a_inst(20);
CPI_A_INST_INTERNAL_20 <= cpi_a_inst(21);
CPI_A_INST_INTERNAL_21 <= cpi_a_inst(22);
CPI_A_INST_INTERNAL_22 <= cpi_a_inst(23);
CPI_A_INST_INTERNAL_23 <= cpi_a_inst(24);
CPI_A_INST_INTERNAL_24 <= cpi_a_inst(25);
CPI_A_INST_INTERNAL_25 <= cpi_a_inst(26);
CPI_A_INST_INTERNAL_26 <= cpi_a_inst(27);
CPI_A_INST_INTERNAL_27 <= cpi_a_inst(28);
CPI_A_INST_INTERNAL_28 <= cpi_a_inst(29);
CPI_A_INST_INTERNAL_29 <= cpi_a_inst(30);
CPI_A_INST_INTERNAL_30 <= cpi_a_inst(31);
CPI_A_CNT_INTERNAL <= cpi_a_cnt(0);
CPI_A_CNT_INTERNAL_0 <= cpi_a_cnt(1);
CPI_A_TRAP_INTERNAL <= cpi_a_trap;
CPI_A_ANNUL_INTERNAL <= cpi_a_annul;
CPI_A_PV_INTERNAL <= cpi_a_pv;
CPI_E_PC_INTERNAL <= cpi_e_pc(0);
CPI_E_PC_INTERNAL_0 <= cpi_e_pc(1);
CPI_E_PC_INTERNAL_1 <= cpi_e_pc(2);
CPI_E_PC_INTERNAL_2 <= cpi_e_pc(3);
CPI_E_PC_INTERNAL_3 <= cpi_e_pc(4);
CPI_E_PC_INTERNAL_4 <= cpi_e_pc(5);
CPI_E_PC_INTERNAL_5 <= cpi_e_pc(6);
CPI_E_PC_INTERNAL_6 <= cpi_e_pc(7);
CPI_E_PC_INTERNAL_7 <= cpi_e_pc(8);
CPI_E_PC_INTERNAL_8 <= cpi_e_pc(9);
CPI_E_PC_INTERNAL_9 <= cpi_e_pc(10);
CPI_E_PC_INTERNAL_10 <= cpi_e_pc(11);
CPI_E_PC_INTERNAL_11 <= cpi_e_pc(12);
CPI_E_PC_INTERNAL_12 <= cpi_e_pc(13);
CPI_E_PC_INTERNAL_13 <= cpi_e_pc(14);
CPI_E_PC_INTERNAL_14 <= cpi_e_pc(15);
CPI_E_PC_INTERNAL_15 <= cpi_e_pc(16);
CPI_E_PC_INTERNAL_16 <= cpi_e_pc(17);
CPI_E_PC_INTERNAL_17 <= cpi_e_pc(18);
CPI_E_PC_INTERNAL_18 <= cpi_e_pc(19);
CPI_E_PC_INTERNAL_19 <= cpi_e_pc(20);
CPI_E_PC_INTERNAL_20 <= cpi_e_pc(21);
CPI_E_PC_INTERNAL_21 <= cpi_e_pc(22);
CPI_E_PC_INTERNAL_22 <= cpi_e_pc(23);
CPI_E_PC_INTERNAL_23 <= cpi_e_pc(24);
CPI_E_PC_INTERNAL_24 <= cpi_e_pc(25);
CPI_E_PC_INTERNAL_25 <= cpi_e_pc(26);
CPI_E_PC_INTERNAL_26 <= cpi_e_pc(27);
CPI_E_PC_INTERNAL_27 <= cpi_e_pc(28);
CPI_E_PC_INTERNAL_28 <= cpi_e_pc(29);
CPI_E_PC_INTERNAL_29 <= cpi_e_pc(30);
CPI_E_PC_INTERNAL_30 <= cpi_e_pc(31);
CPI_E_INST_INTERNAL <= cpi_e_inst(0);
CPI_E_INST_INTERNAL_0 <= cpi_e_inst(1);
CPI_E_INST_INTERNAL_1 <= cpi_e_inst(2);
CPI_E_INST_INTERNAL_2 <= cpi_e_inst(3);
CPI_E_INST_INTERNAL_3 <= cpi_e_inst(4);
CPI_E_INST_INTERNAL_4 <= cpi_e_inst(5);
CPI_E_INST_INTERNAL_5 <= cpi_e_inst(6);
CPI_E_INST_INTERNAL_6 <= cpi_e_inst(7);
CPI_E_INST_INTERNAL_7 <= cpi_e_inst(8);
CPI_E_INST_INTERNAL_8 <= cpi_e_inst(9);
CPI_E_INST_INTERNAL_9 <= cpi_e_inst(10);
CPI_E_INST_INTERNAL_10 <= cpi_e_inst(11);
CPI_E_INST_INTERNAL_11 <= cpi_e_inst(12);
CPI_E_INST_INTERNAL_12 <= cpi_e_inst(13);
CPI_E_INST_INTERNAL_13 <= cpi_e_inst(14);
CPI_E_INST_INTERNAL_14 <= cpi_e_inst(15);
CPI_E_INST_INTERNAL_15 <= cpi_e_inst(16);
CPI_E_INST_INTERNAL_16 <= cpi_e_inst(17);
CPI_E_INST_INTERNAL_17 <= cpi_e_inst(18);
CPI_E_INST_INTERNAL_18 <= cpi_e_inst(19);
CPI_E_INST_INTERNAL_19 <= cpi_e_inst(20);
CPI_E_INST_INTERNAL_20 <= cpi_e_inst(21);
CPI_E_INST_INTERNAL_21 <= cpi_e_inst(22);
CPI_E_INST_INTERNAL_22 <= cpi_e_inst(23);
CPI_E_INST_INTERNAL_23 <= cpi_e_inst(24);
CPI_E_INST_INTERNAL_24 <= cpi_e_inst(25);
CPI_E_INST_INTERNAL_25 <= cpi_e_inst(26);
CPI_E_INST_INTERNAL_26 <= cpi_e_inst(27);
CPI_E_INST_INTERNAL_27 <= cpi_e_inst(28);
CPI_E_INST_INTERNAL_28 <= cpi_e_inst(29);
CPI_E_INST_INTERNAL_29 <= cpi_e_inst(30);
CPI_E_INST_INTERNAL_30 <= cpi_e_inst(31);
CPI_E_CNT_INTERNAL <= cpi_e_cnt(0);
CPI_E_CNT_INTERNAL_0 <= cpi_e_cnt(1);
CPI_E_TRAP_INTERNAL <= cpi_e_trap;
CPI_E_ANNUL_INTERNAL <= cpi_e_annul;
CPI_E_PV_INTERNAL <= cpi_e_pv;
CPI_M_PC_INTERNAL <= cpi_m_pc(0);
CPI_M_PC_INTERNAL_0 <= cpi_m_pc(1);
CPI_M_PC_INTERNAL_1 <= cpi_m_pc(2);
CPI_M_PC_INTERNAL_2 <= cpi_m_pc(3);
CPI_M_PC_INTERNAL_3 <= cpi_m_pc(4);
CPI_M_PC_INTERNAL_4 <= cpi_m_pc(5);
CPI_M_PC_INTERNAL_5 <= cpi_m_pc(6);
CPI_M_PC_INTERNAL_6 <= cpi_m_pc(7);
CPI_M_PC_INTERNAL_7 <= cpi_m_pc(8);
CPI_M_PC_INTERNAL_8 <= cpi_m_pc(9);
CPI_M_PC_INTERNAL_9 <= cpi_m_pc(10);
CPI_M_PC_INTERNAL_10 <= cpi_m_pc(11);
CPI_M_PC_INTERNAL_11 <= cpi_m_pc(12);
CPI_M_PC_INTERNAL_12 <= cpi_m_pc(13);
CPI_M_PC_INTERNAL_13 <= cpi_m_pc(14);
CPI_M_PC_INTERNAL_14 <= cpi_m_pc(15);
CPI_M_PC_INTERNAL_15 <= cpi_m_pc(16);
CPI_M_PC_INTERNAL_16 <= cpi_m_pc(17);
CPI_M_PC_INTERNAL_17 <= cpi_m_pc(18);
CPI_M_PC_INTERNAL_18 <= cpi_m_pc(19);
CPI_M_PC_INTERNAL_19 <= cpi_m_pc(20);
CPI_M_PC_INTERNAL_20 <= cpi_m_pc(21);
CPI_M_PC_INTERNAL_21 <= cpi_m_pc(22);
CPI_M_PC_INTERNAL_22 <= cpi_m_pc(23);
CPI_M_PC_INTERNAL_23 <= cpi_m_pc(24);
CPI_M_PC_INTERNAL_24 <= cpi_m_pc(25);
CPI_M_PC_INTERNAL_25 <= cpi_m_pc(26);
CPI_M_PC_INTERNAL_26 <= cpi_m_pc(27);
CPI_M_PC_INTERNAL_27 <= cpi_m_pc(28);
CPI_M_PC_INTERNAL_28 <= cpi_m_pc(29);
CPI_M_PC_INTERNAL_29 <= cpi_m_pc(30);
CPI_M_PC_INTERNAL_30 <= cpi_m_pc(31);
CPI_M_INST_INTERNAL <= cpi_m_inst(0);
CPI_M_INST_INTERNAL_0 <= cpi_m_inst(1);
CPI_M_INST_INTERNAL_1 <= cpi_m_inst(2);
CPI_M_INST_INTERNAL_2 <= cpi_m_inst(3);
CPI_M_INST_INTERNAL_3 <= cpi_m_inst(4);
CPI_M_INST_INTERNAL_4 <= cpi_m_inst(5);
CPI_M_INST_INTERNAL_5 <= cpi_m_inst(6);
CPI_M_INST_INTERNAL_6 <= cpi_m_inst(7);
CPI_M_INST_INTERNAL_7 <= cpi_m_inst(8);
CPI_M_INST_INTERNAL_8 <= cpi_m_inst(9);
CPI_M_INST_INTERNAL_9 <= cpi_m_inst(10);
CPI_M_INST_INTERNAL_10 <= cpi_m_inst(11);
CPI_M_INST_INTERNAL_11 <= cpi_m_inst(12);
CPI_M_INST_INTERNAL_12 <= cpi_m_inst(13);
CPI_M_INST_INTERNAL_13 <= cpi_m_inst(14);
CPI_M_INST_INTERNAL_14 <= cpi_m_inst(15);
CPI_M_INST_INTERNAL_15 <= cpi_m_inst(16);
CPI_M_INST_INTERNAL_16 <= cpi_m_inst(17);
CPI_M_INST_INTERNAL_17 <= cpi_m_inst(18);
CPI_M_INST_INTERNAL_18 <= cpi_m_inst(19);
CPI_M_INST_INTERNAL_19 <= cpi_m_inst(20);
CPI_M_INST_INTERNAL_20 <= cpi_m_inst(21);
CPI_M_INST_INTERNAL_21 <= cpi_m_inst(22);
CPI_M_INST_INTERNAL_22 <= cpi_m_inst(23);
CPI_M_INST_INTERNAL_23 <= cpi_m_inst(24);
CPI_M_INST_INTERNAL_24 <= cpi_m_inst(25);
CPI_M_INST_INTERNAL_25 <= cpi_m_inst(26);
CPI_M_INST_INTERNAL_26 <= cpi_m_inst(27);
CPI_M_INST_INTERNAL_27 <= cpi_m_inst(28);
CPI_M_INST_INTERNAL_28 <= cpi_m_inst(29);
CPI_M_INST_INTERNAL_29 <= cpi_m_inst(30);
CPI_M_INST_INTERNAL_30 <= cpi_m_inst(31);
CPI_M_CNT_INTERNAL <= cpi_m_cnt(0);
CPI_M_CNT_INTERNAL_0 <= cpi_m_cnt(1);
CPI_M_TRAP_INTERNAL <= cpi_m_trap;
CPI_M_ANNUL_INTERNAL <= cpi_m_annul;
CPI_M_PV_INTERNAL <= cpi_m_pv;
CPI_X_PC_INTERNAL <= cpi_x_pc(0);
CPI_X_PC_INTERNAL_0 <= cpi_x_pc(1);
CPI_X_PC_INTERNAL_1 <= cpi_x_pc(2);
CPI_X_PC_INTERNAL_2 <= cpi_x_pc(3);
CPI_X_PC_INTERNAL_3 <= cpi_x_pc(4);
CPI_X_PC_INTERNAL_4 <= cpi_x_pc(5);
CPI_X_PC_INTERNAL_5 <= cpi_x_pc(6);
CPI_X_PC_INTERNAL_6 <= cpi_x_pc(7);
CPI_X_PC_INTERNAL_7 <= cpi_x_pc(8);
CPI_X_PC_INTERNAL_8 <= cpi_x_pc(9);
CPI_X_PC_INTERNAL_9 <= cpi_x_pc(10);
CPI_X_PC_INTERNAL_10 <= cpi_x_pc(11);
CPI_X_PC_INTERNAL_11 <= cpi_x_pc(12);
CPI_X_PC_INTERNAL_12 <= cpi_x_pc(13);
CPI_X_PC_INTERNAL_13 <= cpi_x_pc(14);
CPI_X_PC_INTERNAL_14 <= cpi_x_pc(15);
CPI_X_PC_INTERNAL_15 <= cpi_x_pc(16);
CPI_X_PC_INTERNAL_16 <= cpi_x_pc(17);
CPI_X_PC_INTERNAL_17 <= cpi_x_pc(18);
CPI_X_PC_INTERNAL_18 <= cpi_x_pc(19);
CPI_X_PC_INTERNAL_19 <= cpi_x_pc(20);
CPI_X_PC_INTERNAL_20 <= cpi_x_pc(21);
CPI_X_PC_INTERNAL_21 <= cpi_x_pc(22);
CPI_X_PC_INTERNAL_22 <= cpi_x_pc(23);
CPI_X_PC_INTERNAL_23 <= cpi_x_pc(24);
CPI_X_PC_INTERNAL_24 <= cpi_x_pc(25);
CPI_X_PC_INTERNAL_25 <= cpi_x_pc(26);
CPI_X_PC_INTERNAL_26 <= cpi_x_pc(27);
CPI_X_PC_INTERNAL_27 <= cpi_x_pc(28);
CPI_X_PC_INTERNAL_28 <= cpi_x_pc(29);
CPI_X_PC_INTERNAL_29 <= cpi_x_pc(30);
CPI_X_PC_INTERNAL_30 <= cpi_x_pc(31);
CPI_X_INST_INTERNAL <= cpi_x_inst(0);
CPI_X_INST_INTERNAL_0 <= cpi_x_inst(1);
CPI_X_INST_INTERNAL_1 <= cpi_x_inst(2);
CPI_X_INST_INTERNAL_2 <= cpi_x_inst(3);
CPI_X_INST_INTERNAL_3 <= cpi_x_inst(4);
CPI_X_INST_INTERNAL_4 <= cpi_x_inst(5);
CPI_X_INST_INTERNAL_5 <= cpi_x_inst(6);
CPI_X_INST_INTERNAL_6 <= cpi_x_inst(7);
CPI_X_INST_INTERNAL_7 <= cpi_x_inst(8);
CPI_X_INST_INTERNAL_8 <= cpi_x_inst(9);
CPI_X_INST_INTERNAL_9 <= cpi_x_inst(10);
CPI_X_INST_INTERNAL_10 <= cpi_x_inst(11);
CPI_X_INST_INTERNAL_11 <= cpi_x_inst(12);
CPI_X_INST_INTERNAL_12 <= cpi_x_inst(13);
CPI_X_INST_INTERNAL_13 <= cpi_x_inst(14);
CPI_X_INST_INTERNAL_14 <= cpi_x_inst(15);
CPI_X_INST_INTERNAL_15 <= cpi_x_inst(16);
CPI_X_INST_INTERNAL_16 <= cpi_x_inst(17);
CPI_X_INST_INTERNAL_17 <= cpi_x_inst(18);
CPI_X_INST_INTERNAL_18 <= cpi_x_inst(19);
CPI_X_INST_INTERNAL_19 <= cpi_x_inst(20);
CPI_X_INST_INTERNAL_20 <= cpi_x_inst(21);
CPI_X_INST_INTERNAL_21 <= cpi_x_inst(22);
CPI_X_INST_INTERNAL_22 <= cpi_x_inst(23);
CPI_X_INST_INTERNAL_23 <= cpi_x_inst(24);
CPI_X_INST_INTERNAL_24 <= cpi_x_inst(25);
CPI_X_INST_INTERNAL_25 <= cpi_x_inst(26);
CPI_X_INST_INTERNAL_26 <= cpi_x_inst(27);
CPI_X_INST_INTERNAL_27 <= cpi_x_inst(28);
CPI_X_INST_INTERNAL_28 <= cpi_x_inst(29);
CPI_X_INST_INTERNAL_29 <= cpi_x_inst(30);
CPI_X_INST_INTERNAL_30 <= cpi_x_inst(31);
CPI_X_CNT_INTERNAL <= cpi_x_cnt(0);
CPI_X_CNT_INTERNAL_0 <= cpi_x_cnt(1);
CPI_X_TRAP_INTERNAL <= cpi_x_trap;
CPI_X_ANNUL_INTERNAL <= cpi_x_annul;
CPI_X_PV_INTERNAL <= cpi_x_pv;
CPI_LDDATA_INTERNAL <= cpi_lddata(0);
CPI_LDDATA_INTERNAL_0 <= cpi_lddata(1);
CPI_LDDATA_INTERNAL_1 <= cpi_lddata(2);
CPI_LDDATA_INTERNAL_2 <= cpi_lddata(3);
CPI_LDDATA_INTERNAL_3 <= cpi_lddata(4);
CPI_LDDATA_INTERNAL_4 <= cpi_lddata(5);
CPI_LDDATA_INTERNAL_5 <= cpi_lddata(6);
CPI_LDDATA_INTERNAL_6 <= cpi_lddata(7);
CPI_LDDATA_INTERNAL_7 <= cpi_lddata(8);
CPI_LDDATA_INTERNAL_8 <= cpi_lddata(9);
CPI_LDDATA_INTERNAL_9 <= cpi_lddata(10);
CPI_LDDATA_INTERNAL_10 <= cpi_lddata(11);
CPI_LDDATA_INTERNAL_11 <= cpi_lddata(12);
CPI_LDDATA_INTERNAL_12 <= cpi_lddata(13);
CPI_LDDATA_INTERNAL_13 <= cpi_lddata(14);
CPI_LDDATA_INTERNAL_14 <= cpi_lddata(15);
CPI_LDDATA_INTERNAL_15 <= cpi_lddata(16);
CPI_LDDATA_INTERNAL_16 <= cpi_lddata(17);
CPI_LDDATA_INTERNAL_17 <= cpi_lddata(18);
CPI_LDDATA_INTERNAL_18 <= cpi_lddata(19);
CPI_LDDATA_INTERNAL_19 <= cpi_lddata(20);
CPI_LDDATA_INTERNAL_20 <= cpi_lddata(21);
CPI_LDDATA_INTERNAL_21 <= cpi_lddata(22);
CPI_LDDATA_INTERNAL_22 <= cpi_lddata(23);
CPI_LDDATA_INTERNAL_23 <= cpi_lddata(24);
CPI_LDDATA_INTERNAL_24 <= cpi_lddata(25);
CPI_LDDATA_INTERNAL_25 <= cpi_lddata(26);
CPI_LDDATA_INTERNAL_26 <= cpi_lddata(27);
CPI_LDDATA_INTERNAL_27 <= cpi_lddata(28);
CPI_LDDATA_INTERNAL_28 <= cpi_lddata(29);
CPI_LDDATA_INTERNAL_29 <= cpi_lddata(30);
CPI_LDDATA_INTERNAL_30 <= cpi_lddata(31);
CPI_DBG_ENABLE_INTERNAL <= cpi_dbg_enable;
CPI_DBG_WRITE_INTERNAL <= cpi_dbg_write;
CPI_DBG_FSR_INTERNAL <= cpi_dbg_fsr;
CPI_DBG_ADDR_INTERNAL <= cpi_dbg_addr(0);
CPI_DBG_ADDR_INTERNAL_0 <= cpi_dbg_addr(1);
CPI_DBG_ADDR_INTERNAL_1 <= cpi_dbg_addr(2);
CPI_DBG_ADDR_INTERNAL_2 <= cpi_dbg_addr(3);
CPI_DBG_ADDR_INTERNAL_3 <= cpi_dbg_addr(4);
CPI_DBG_DATA_INTERNAL <= cpi_dbg_data(0);
CPI_DBG_DATA_INTERNAL_0 <= cpi_dbg_data(1);
CPI_DBG_DATA_INTERNAL_1 <= cpi_dbg_data(2);
CPI_DBG_DATA_INTERNAL_2 <= cpi_dbg_data(3);
CPI_DBG_DATA_INTERNAL_3 <= cpi_dbg_data(4);
CPI_DBG_DATA_INTERNAL_4 <= cpi_dbg_data(5);
CPI_DBG_DATA_INTERNAL_5 <= cpi_dbg_data(6);
CPI_DBG_DATA_INTERNAL_6 <= cpi_dbg_data(7);
CPI_DBG_DATA_INTERNAL_7 <= cpi_dbg_data(8);
CPI_DBG_DATA_INTERNAL_8 <= cpi_dbg_data(9);
CPI_DBG_DATA_INTERNAL_9 <= cpi_dbg_data(10);
CPI_DBG_DATA_INTERNAL_10 <= cpi_dbg_data(11);
CPI_DBG_DATA_INTERNAL_11 <= cpi_dbg_data(12);
CPI_DBG_DATA_INTERNAL_12 <= cpi_dbg_data(13);
CPI_DBG_DATA_INTERNAL_13 <= cpi_dbg_data(14);
CPI_DBG_DATA_INTERNAL_14 <= cpi_dbg_data(15);
CPI_DBG_DATA_INTERNAL_15 <= cpi_dbg_data(16);
CPI_DBG_DATA_INTERNAL_16 <= cpi_dbg_data(17);
CPI_DBG_DATA_INTERNAL_17 <= cpi_dbg_data(18);
CPI_DBG_DATA_INTERNAL_18 <= cpi_dbg_data(19);
CPI_DBG_DATA_INTERNAL_19 <= cpi_dbg_data(20);
CPI_DBG_DATA_INTERNAL_20 <= cpi_dbg_data(21);
CPI_DBG_DATA_INTERNAL_21 <= cpi_dbg_data(22);
CPI_DBG_DATA_INTERNAL_22 <= cpi_dbg_data(23);
CPI_DBG_DATA_INTERNAL_23 <= cpi_dbg_data(24);
CPI_DBG_DATA_INTERNAL_24 <= cpi_dbg_data(25);
CPI_DBG_DATA_INTERNAL_25 <= cpi_dbg_data(26);
CPI_DBG_DATA_INTERNAL_26 <= cpi_dbg_data(27);
CPI_DBG_DATA_INTERNAL_27 <= cpi_dbg_data(28);
CPI_DBG_DATA_INTERNAL_28 <= cpi_dbg_data(29);
CPI_DBG_DATA_INTERNAL_29 <= cpi_dbg_data(30);
CPI_DBG_DATA_INTERNAL_30 <= cpi_dbg_data(31);
RFO1_DATA1_INTERNAL <= rfo1_data1(0);
RFO1_DATA1_INTERNAL_0 <= rfo1_data1(1);
RFO1_DATA1_INTERNAL_1 <= rfo1_data1(2);
RFO1_DATA1_INTERNAL_2 <= rfo1_data1(3);
RFO1_DATA1_INTERNAL_3 <= rfo1_data1(4);
RFO1_DATA1_INTERNAL_4 <= rfo1_data1(5);
RFO1_DATA1_INTERNAL_5 <= rfo1_data1(6);
RFO1_DATA1_INTERNAL_6 <= rfo1_data1(7);
RFO1_DATA1_INTERNAL_7 <= rfo1_data1(8);
RFO1_DATA1_INTERNAL_8 <= rfo1_data1(9);
RFO1_DATA1_INTERNAL_9 <= rfo1_data1(10);
RFO1_DATA1_INTERNAL_10 <= rfo1_data1(11);
RFO1_DATA1_INTERNAL_11 <= rfo1_data1(12);
RFO1_DATA1_INTERNAL_12 <= rfo1_data1(13);
RFO1_DATA1_INTERNAL_13 <= rfo1_data1(14);
RFO1_DATA1_INTERNAL_14 <= rfo1_data1(15);
RFO1_DATA1_INTERNAL_15 <= rfo1_data1(16);
RFO1_DATA1_INTERNAL_16 <= rfo1_data1(17);
RFO1_DATA1_INTERNAL_17 <= rfo1_data1(18);
RFO1_DATA1_INTERNAL_18 <= rfo1_data1(19);
RFO1_DATA1_INTERNAL_19 <= rfo1_data1(20);
RFO1_DATA1_INTERNAL_20 <= rfo1_data1(21);
RFO1_DATA1_INTERNAL_21 <= rfo1_data1(22);
RFO1_DATA1_INTERNAL_22 <= rfo1_data1(23);
RFO1_DATA1_INTERNAL_23 <= rfo1_data1(24);
RFO1_DATA1_INTERNAL_24 <= rfo1_data1(25);
RFO1_DATA1_INTERNAL_25 <= rfo1_data1(26);
RFO1_DATA1_INTERNAL_26 <= rfo1_data1(27);
RFO1_DATA1_INTERNAL_27 <= rfo1_data1(28);
RFO1_DATA1_INTERNAL_28 <= rfo1_data1(29);
RFO1_DATA1_INTERNAL_29 <= rfo1_data1(30);
RFO1_DATA1_INTERNAL_30 <= rfo1_data1(31);
RFO1_DATA2_INTERNAL <= rfo1_data2(0);
RFO1_DATA2_INTERNAL_0 <= rfo1_data2(1);
RFO1_DATA2_INTERNAL_1 <= rfo1_data2(2);
RFO1_DATA2_INTERNAL_2 <= rfo1_data2(3);
RFO1_DATA2_INTERNAL_3 <= rfo1_data2(4);
RFO1_DATA2_INTERNAL_4 <= rfo1_data2(5);
RFO1_DATA2_INTERNAL_5 <= rfo1_data2(6);
RFO1_DATA2_INTERNAL_6 <= rfo1_data2(7);
RFO1_DATA2_INTERNAL_7 <= rfo1_data2(8);
RFO1_DATA2_INTERNAL_8 <= rfo1_data2(9);
RFO1_DATA2_INTERNAL_9 <= rfo1_data2(10);
RFO1_DATA2_INTERNAL_10 <= rfo1_data2(11);
RFO1_DATA2_INTERNAL_11 <= rfo1_data2(12);
RFO1_DATA2_INTERNAL_12 <= rfo1_data2(13);
RFO1_DATA2_INTERNAL_13 <= rfo1_data2(14);
RFO1_DATA2_INTERNAL_14 <= rfo1_data2(15);
RFO1_DATA2_INTERNAL_15 <= rfo1_data2(16);
RFO1_DATA2_INTERNAL_16 <= rfo1_data2(17);
RFO1_DATA2_INTERNAL_17 <= rfo1_data2(18);
RFO1_DATA2_INTERNAL_18 <= rfo1_data2(19);
RFO1_DATA2_INTERNAL_19 <= rfo1_data2(20);
RFO1_DATA2_INTERNAL_20 <= rfo1_data2(21);
RFO1_DATA2_INTERNAL_21 <= rfo1_data2(22);
RFO1_DATA2_INTERNAL_22 <= rfo1_data2(23);
RFO1_DATA2_INTERNAL_23 <= rfo1_data2(24);
RFO1_DATA2_INTERNAL_24 <= rfo1_data2(25);
RFO1_DATA2_INTERNAL_25 <= rfo1_data2(26);
RFO1_DATA2_INTERNAL_26 <= rfo1_data2(27);
RFO1_DATA2_INTERNAL_27 <= rfo1_data2(28);
RFO1_DATA2_INTERNAL_28 <= rfo1_data2(29);
RFO1_DATA2_INTERNAL_29 <= rfo1_data2(30);
RFO1_DATA2_INTERNAL_30 <= rfo1_data2(31);
RFO2_DATA1_INTERNAL <= rfo2_data1(0);
RFO2_DATA1_INTERNAL_0 <= rfo2_data1(1);
RFO2_DATA1_INTERNAL_1 <= rfo2_data1(2);
RFO2_DATA1_INTERNAL_2 <= rfo2_data1(3);
RFO2_DATA1_INTERNAL_3 <= rfo2_data1(4);
RFO2_DATA1_INTERNAL_4 <= rfo2_data1(5);
RFO2_DATA1_INTERNAL_5 <= rfo2_data1(6);
RFO2_DATA1_INTERNAL_6 <= rfo2_data1(7);
RFO2_DATA1_INTERNAL_7 <= rfo2_data1(8);
RFO2_DATA1_INTERNAL_8 <= rfo2_data1(9);
RFO2_DATA1_INTERNAL_9 <= rfo2_data1(10);
RFO2_DATA1_INTERNAL_10 <= rfo2_data1(11);
RFO2_DATA1_INTERNAL_11 <= rfo2_data1(12);
RFO2_DATA1_INTERNAL_12 <= rfo2_data1(13);
RFO2_DATA1_INTERNAL_13 <= rfo2_data1(14);
RFO2_DATA1_INTERNAL_14 <= rfo2_data1(15);
RFO2_DATA1_INTERNAL_15 <= rfo2_data1(16);
RFO2_DATA1_INTERNAL_16 <= rfo2_data1(17);
RFO2_DATA1_INTERNAL_17 <= rfo2_data1(18);
RFO2_DATA1_INTERNAL_18 <= rfo2_data1(19);
RFO2_DATA1_INTERNAL_19 <= rfo2_data1(20);
RFO2_DATA1_INTERNAL_20 <= rfo2_data1(21);
RFO2_DATA1_INTERNAL_21 <= rfo2_data1(22);
RFO2_DATA1_INTERNAL_22 <= rfo2_data1(23);
RFO2_DATA1_INTERNAL_23 <= rfo2_data1(24);
RFO2_DATA1_INTERNAL_24 <= rfo2_data1(25);
RFO2_DATA1_INTERNAL_25 <= rfo2_data1(26);
RFO2_DATA1_INTERNAL_26 <= rfo2_data1(27);
RFO2_DATA1_INTERNAL_27 <= rfo2_data1(28);
RFO2_DATA1_INTERNAL_28 <= rfo2_data1(29);
RFO2_DATA1_INTERNAL_29 <= rfo2_data1(30);
RFO2_DATA1_INTERNAL_30 <= rfo2_data1(31);
RFO2_DATA2_INTERNAL <= rfo2_data2(0);
RFO2_DATA2_INTERNAL_0 <= rfo2_data2(1);
RFO2_DATA2_INTERNAL_1 <= rfo2_data2(2);
RFO2_DATA2_INTERNAL_2 <= rfo2_data2(3);
RFO2_DATA2_INTERNAL_3 <= rfo2_data2(4);
RFO2_DATA2_INTERNAL_4 <= rfo2_data2(5);
RFO2_DATA2_INTERNAL_5 <= rfo2_data2(6);
RFO2_DATA2_INTERNAL_6 <= rfo2_data2(7);
RFO2_DATA2_INTERNAL_7 <= rfo2_data2(8);
RFO2_DATA2_INTERNAL_8 <= rfo2_data2(9);
RFO2_DATA2_INTERNAL_9 <= rfo2_data2(10);
RFO2_DATA2_INTERNAL_10 <= rfo2_data2(11);
RFO2_DATA2_INTERNAL_11 <= rfo2_data2(12);
RFO2_DATA2_INTERNAL_12 <= rfo2_data2(13);
RFO2_DATA2_INTERNAL_13 <= rfo2_data2(14);
RFO2_DATA2_INTERNAL_14 <= rfo2_data2(15);
RFO2_DATA2_INTERNAL_15 <= rfo2_data2(16);
RFO2_DATA2_INTERNAL_16 <= rfo2_data2(17);
RFO2_DATA2_INTERNAL_17 <= rfo2_data2(18);
RFO2_DATA2_INTERNAL_18 <= rfo2_data2(19);
RFO2_DATA2_INTERNAL_19 <= rfo2_data2(20);
RFO2_DATA2_INTERNAL_20 <= rfo2_data2(21);
RFO2_DATA2_INTERNAL_21 <= rfo2_data2(22);
RFO2_DATA2_INTERNAL_22 <= rfo2_data2(23);
RFO2_DATA2_INTERNAL_23 <= rfo2_data2(24);
RFO2_DATA2_INTERNAL_24 <= rfo2_data2(25);
RFO2_DATA2_INTERNAL_25 <= rfo2_data2(26);
RFO2_DATA2_INTERNAL_26 <= rfo2_data2(27);
RFO2_DATA2_INTERNAL_27 <= rfo2_data2(28);
RFO2_DATA2_INTERNAL_28 <= rfo2_data2(29);
RFO2_DATA2_INTERNAL_29 <= rfo2_data2(30);
RFO2_DATA2_INTERNAL_30 <= rfo2_data2(31);
end beh;

