------------------------------------------------------------------------------
--  This file is a part of the GRLIB VHDL IP LIBRARY
--  Copyright (C) 2006-2010, Aeroflex Gaisler AB - all rights reserved.
--
-- ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN 
-- ACCORDANCE WITH THE GAISLER LICENSE AGREEMENT AND MUST BE APPROVED 
-- IN ADVANCE IN WRITING. 
-----------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
library UNISIM;
use UNISIM.vcomponents.all;
use UNISIM.all;

entity grlfpw_0_unisim is
port(
  rst :  in std_logic;
  clk :  in std_logic;
  holdn :  in std_logic;
  cpi_flush :  in std_logic;
  cpi_exack :  in std_logic;
  cpi_a_rs1 : in std_logic_vector (4 downto 0);
  cpi_d_pc : in std_logic_vector (31 downto 0);
  cpi_d_inst : in std_logic_vector (31 downto 0);
  cpi_d_cnt : in std_logic_vector (1 downto 0);
  cpi_d_trap :  in std_logic;
  cpi_d_annul :  in std_logic;
  cpi_d_pv :  in std_logic;
  cpi_a_pc : in std_logic_vector (31 downto 0);
  cpi_a_inst : in std_logic_vector (31 downto 0);
  cpi_a_cnt : in std_logic_vector (1 downto 0);
  cpi_a_trap :  in std_logic;
  cpi_a_annul :  in std_logic;
  cpi_a_pv :  in std_logic;
  cpi_e_pc : in std_logic_vector (31 downto 0);
  cpi_e_inst : in std_logic_vector (31 downto 0);
  cpi_e_cnt : in std_logic_vector (1 downto 0);
  cpi_e_trap :  in std_logic;
  cpi_e_annul :  in std_logic;
  cpi_e_pv :  in std_logic;
  cpi_m_pc : in std_logic_vector (31 downto 0);
  cpi_m_inst : in std_logic_vector (31 downto 0);
  cpi_m_cnt : in std_logic_vector (1 downto 0);
  cpi_m_trap :  in std_logic;
  cpi_m_annul :  in std_logic;
  cpi_m_pv :  in std_logic;
  cpi_x_pc : in std_logic_vector (31 downto 0);
  cpi_x_inst : in std_logic_vector (31 downto 0);
  cpi_x_cnt : in std_logic_vector (1 downto 0);
  cpi_x_trap :  in std_logic;
  cpi_x_annul :  in std_logic;
  cpi_x_pv :  in std_logic;
  cpi_lddata : in std_logic_vector (31 downto 0);
  cpi_dbg_enable :  in std_logic;
  cpi_dbg_write :  in std_logic;
  cpi_dbg_fsr :  in std_logic;
  cpi_dbg_addr : in std_logic_vector (4 downto 0);
  cpi_dbg_data : in std_logic_vector (31 downto 0);
  cpo_data : out std_logic_vector (31 downto 0);
  cpo_exc :  out std_logic;
  cpo_cc : out std_logic_vector (1 downto 0);
  cpo_ccv :  out std_logic;
  cpo_ldlock :  out std_logic;
  cpo_holdn :  out std_logic;
  cpo_dbg_data : out std_logic_vector (31 downto 0);
  rfi1_rd1addr : out std_logic_vector (3 downto 0);
  rfi1_rd2addr : out std_logic_vector (3 downto 0);
  rfi1_wraddr : out std_logic_vector (3 downto 0);
  rfi1_wrdata : out std_logic_vector (31 downto 0);
  rfi1_ren1 :  out std_logic;
  rfi1_ren2 :  out std_logic;
  rfi1_wren :  out std_logic;
  rfi2_rd1addr : out std_logic_vector (3 downto 0);
  rfi2_rd2addr : out std_logic_vector (3 downto 0);
  rfi2_wraddr : out std_logic_vector (3 downto 0);
  rfi2_wrdata : out std_logic_vector (31 downto 0);
  rfi2_ren1 :  out std_logic;
  rfi2_ren2 :  out std_logic;
  rfi2_wren :  out std_logic;
  rfo1_data1 : in std_logic_vector (31 downto 0);
  rfo1_data2 : in std_logic_vector (31 downto 0);
  rfo2_data1 : in std_logic_vector (31 downto 0);
  rfo2_data2 : in std_logic_vector (31 downto 0));
end grlfpw_0_unisim;

architecture beh of grlfpw_0_unisim is
  component FDRSE
	generic ( INIT : bit := '0');
	port (  Q : out std_ulogic;
		C : in std_ulogic;
		CE : in std_ulogic;
		D : in std_ulogic;
		R : in std_ulogic;
		S : in std_ulogic);
  end component;

  component FDR
	generic ( INIT : bit := '0');
	port (  Q : out std_ulogic;
		C : in std_ulogic;
		D : in std_ulogic;
		R : in std_ulogic);
  end component;

  component FDRE
	generic ( INIT : bit := '0');
	port (  Q : out std_ulogic;
		C : in std_ulogic;
		CE : in std_ulogic;
		D : in std_ulogic;
		R : in std_ulogic);
  end component;

  component FD
	generic ( INIT : bit := '0');
	port (  Q : out std_ulogic;
		C : in std_ulogic;
		D : in std_ulogic);
  end component;

  component FDRS
	generic ( INIT : bit := '0');
	port (  Q : out std_ulogic;
		C : in std_ulogic;
		D : in std_ulogic;
		R : in std_ulogic;
		S : in std_ulogic);
  end component;

  component FDE
	generic ( INIT : bit := '0');
	port (  Q : out std_ulogic;
		C : in std_ulogic;
		CE : in std_ulogic;
		D : in std_ulogic);
  end component;

  component MUXF5
	port (  O : out std_ulogic;
		I0 : in std_ulogic;
		I1 : in std_ulogic;
		S : in std_ulogic);
  end component;

  component VCC
	port ( P : out std_ulogic := '1');
  end component;

  component GND
	port ( G : out std_ulogic := '0');
  end component;

component INV
	port
	(
		O : out std_ulogic;
		I : in std_ulogic
	);
end component;
component LUT2_L
	generic
	(
		INIT : bit_vector := X"0"
	);
	port
	(
		LO : out std_ulogic;
		I0 : in std_ulogic;
		I1 : in std_ulogic
	);
end component;
component LUT4
	generic
	(
		INIT : bit_vector := X"0000"
	);
	port
	(
		O : out std_ulogic;
		I0 : in std_ulogic;
		I1 : in std_ulogic;
		I2 : in std_ulogic;
		I3 : in std_ulogic
	);
end component;
component LUT3
	generic
	(
		INIT : bit_vector := X"00"
	);
	port
	(
		O : out std_ulogic;
		I0 : in std_ulogic;
		I1 : in std_ulogic;
		I2 : in std_ulogic
	);
end component;
component LUT2
	generic
	(
		INIT : bit_vector := X"0"
	);
	port
	(
		O : out std_ulogic;
		I0 : in std_ulogic;
		I1 : in std_ulogic
	);
end component;
component FDC
	generic
	(
		INIT : bit := '0'
	);
	port
	(
		Q : out std_ulogic;
		C : in std_ulogic;
		CLR : in std_ulogic;
		D : in std_ulogic
	);
end component;
component LUT3_L
	generic
	(
		INIT : bit_vector := X"00"
	);
	port
	(
		LO : out std_ulogic;
		I0 : in std_ulogic;
		I1 : in std_ulogic;
		I2 : in std_ulogic
	);
end component;
component LUT1
	generic
	(
		INIT : bit_vector := X"0"
	);
	port
	(
		O : out std_ulogic;
		I0 : in std_ulogic
	);
end component;
component LUT4_L
	generic
	(
		INIT : bit_vector := X"0000"
	);
	port
	(
		LO : out std_ulogic;
		I0 : in std_ulogic;
		I1 : in std_ulogic;
		I2 : in std_ulogic;
		I3 : in std_ulogic
	);
end component;
component FDCE
	generic
	(
		INIT : bit := '0'
	);
	port
	(
		Q : out std_ulogic;
		C : in std_ulogic;
		CE : in std_ulogic;
		CLR : in std_ulogic;
		D : in std_ulogic
	);
end component;
component FDC_1
	generic
	(
		INIT : bit := '0'
	);
	port
	(
		Q : out std_ulogic;
		C : in std_ulogic;
		CLR : in std_ulogic;
		D : in std_ulogic
	);
end component;
component FDP
	generic
	(
		INIT : bit := '1'
	);
	port
	(
		Q : out std_ulogic;
		C : in std_ulogic;
		D : in std_ulogic;
		PRE : in std_ulogic
	);
end component;
component FDS
	generic
	(
		INIT : bit := '1'
	);
	port
	(
		Q : out std_ulogic;
		C : in std_ulogic;
		D : in std_ulogic;
		S : in std_ulogic
	);
end component;
component MUXCY
	port
	(
		O : out std_ulogic;
		CI : in std_ulogic;
		DI : in std_ulogic;
		S : in std_ulogic
	);
end component;
component LUT1_L
	generic
	(
		INIT : bit_vector := X"0"
	);
	port
	(
		LO : out std_ulogic;
		I0 : in std_ulogic
	);
end component;
component MUXF6
	port
	(
		O : out std_ulogic;
		I0 : in std_ulogic;
		I1 : in std_ulogic;
		S : in std_ulogic
	);
end component;
component MUXF5_D
	port
	(
		LO : out std_ulogic;
		O : out std_ulogic;
		I0 : in std_ulogic;
		I1 : in std_ulogic;
		S : in std_ulogic
	);
end component;
component XORCY
	port
	(
		O : out std_ulogic;
		CI : in std_ulogic;
		LI : in std_ulogic
	);
end component;
component MUXCY_L
	port
	(
		LO : out std_ulogic;
		CI : in std_ulogic;
		DI : in std_ulogic;
		S : in std_ulogic
	);
end component;
component FDSE
	generic
	(
		INIT : bit := '1'
	);
	port
	(
		Q : out std_ulogic;
		C : in std_ulogic;
		CE : in std_ulogic;
		D : in std_ulogic;
		S : in std_ulogic
	);
end component;
component MULT_AND
	port
	(
		LO : out std_ulogic;
		I0 : in std_ulogic;
		I1 : in std_ulogic
	);
end component;

component SRL16E
	generic
	(
		INIT : bit_vector := X"0000"
	);
	port
	(
		Q : out STD_ULOGIC;
		A0 : in STD_ULOGIC;
		A1 : in STD_ULOGIC;
		A2 : in STD_ULOGIC;
		A3 : in STD_ULOGIC;
		CE : in STD_ULOGIC;
		CLK : in STD_ULOGIC;
		D : in STD_ULOGIC
	);
end component;

  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL : std_logic_vector (16 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_5 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_4 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_13 : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_14 : std_logic_vector (4 to 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_16 : std_logic_vector (6 to 6);
  signal CPI_D_INST_I : std_logic_vector (31 downto 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_1_I : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_I : std_logic_vector (43 downto 15);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_RESVEC : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL : std_logic_vector (85 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_18 : std_logic_vector (74 to 74);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14 : std_logic_vector (77 to 77);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT : std_logic_vector (7 downto 0);
  signal GRLFPC2_0_R_I_EXC : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_FPO_EXC : std_logic_vector (3 downto 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH : std_logic_vector (377 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE : std_logic_vector (12 downto 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS : std_logic_vector (9 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_MIXOIN : std_logic_vector (0 to 0);
  signal GRLFPC2_0_FPO_EXP : std_logic_vector (10 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS : std_logic_vector (55 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN4_TEMP : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0 : std_logic_vector (57 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1 : std_logic_vector (57 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_I : std_logic_vector (375 to 375);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_I : std_logic_vector (375 to 375);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0 : std_logic_vector (173 downto 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14_M : std_logic_vector (171 downto 142);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M : std_logic_vector (174 downto 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M : std_logic_vector (47 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0_M : std_logic_vector (1 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M : std_logic_vector (57 downto 42);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0_I_M : std_logic_vector (55 to 55);
  signal GRLFPC2_0_R_A_RS2 : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG : std_logic_vector (7 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPYBUS_2 : std_logic_vector (6 to 6);
  signal GRLFPC2_0_R_STATE : std_logic_vector (1 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3 : std_logic_vector (55 downto 0);
  signal GRLFPC2_0_R_FSR_TEM : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_COMB_MEXC_1 : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_LIB : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2 : std_logic_vector (30 downto 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_CONDITIONAL : std_logic_vector (6 to 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN : std_logic_vector (8 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive : std_logic_vector (8 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_1 : std_logic_vector (12 downto 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_FAST : std_logic_vector (17 downto 16);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS : std_logic_vector (57 downto 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_T_3_I_A2_0_0 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_4 : std_logic_vector (6 downto 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_5 : std_logic_vector (6 downto 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_DREG_FAST : std_logic_vector (53 downto 51);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_FAST : std_logic_vector (376 downto 375);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1 : std_logic_vector (3 downto 0);
  signal GRLFPC2_0_R_A_RS1 : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_R_FSR_CEXC : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_R_FSR_AEXC : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_R_FSR_RD : std_logic_vector (1 downto 0);
  signal GRLFPC2_0_R_FSR_FTT : std_logic_vector (2 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4 : std_logic_vector (57 downto 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M2 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_2 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23 : std_logic_vector (113 to 113);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_1 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_R_I_INST : std_logic_vector (31 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1 : std_logic_vector (51 to 51);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_EXPBREGLC_1 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8 : std_logic_vector (57 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14_M_0 : std_logic_vector (171 to 171);
  signal GRLFPC2_0_COMB_V_FSR_RD_1_M1 : std_logic_vector (1 downto 0);
  signal GRLFPC2_0_COMB_V_FSR_TEM_1_M1 : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_COMB_V_FSR_FCC_1_M0 : std_logic_vector (1 downto 0);
  signal GRLFPC2_0_OP1 : std_logic_vector (63 downto 32);
  signal GRLFPC2_0_OP2 : std_logic_vector (63 downto 32);
  signal GRLFPC2_0_R_I_RES : std_logic_vector (63 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_114_1_1_0 : std_logic_vector (56 to 56);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M13 : std_logic_vector (2 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M12 : std_logic_vector (2 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_1 : std_logic_vector (68 to 68);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1 : std_logic_vector (4 downto 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_2_1 : std_logic_vector (1 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2 : std_logic_vector (56 downto 1);
  signal GRLFPC2_0_COMB_WRADDR_5 : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_1 : std_logic_vector (54 downto 0);
  signal GRLFPC2_0_COMB_RS2_1 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1 : std_logic_vector (25 downto 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19 : std_logic_vector (83 downto 61);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M14 : std_logic_vector (3 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_62_1 : std_logic_vector (51 to 51);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_50 : std_logic_vector (7 to 7);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_6 : std_logic_vector (51 to 51);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_49 : std_logic_vector (8 to 8);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_43 : std_logic_vector (14 to 14);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_36 : std_logic_vector (21 to 21);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_31 : std_logic_vector (26 to 26);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_39 : std_logic_vector (18 to 18);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_27 : std_logic_vector (30 to 30);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_32 : std_logic_vector (25 to 25);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_23 : std_logic_vector (34 to 34);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_28 : std_logic_vector (29 to 29);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_16 : std_logic_vector (41 to 41);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_18 : std_logic_vector (39 to 39);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_20 : std_logic_vector (37 to 37);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_25 : std_logic_vector (32 to 32);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_46 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_17 : std_logic_vector (40 to 40);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_37 : std_logic_vector (20 to 20);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_29 : std_logic_vector (28 to 28);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_113_0 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SBLSBS_1_0 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_11 : std_logic_vector (46 to 46);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_22 : std_logic_vector (35 to 35);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_45 : std_logic_vector (12 to 12);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_42 : std_logic_vector (15 to 15);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_40 : std_logic_vector (17 to 17);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_53 : std_logic_vector (4 to 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_26 : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_12 : std_logic_vector (45 to 45);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_48 : std_logic_vector (9 to 9);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_51 : std_logic_vector (6 to 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_15 : std_logic_vector (42 to 42);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SBLSBS_0 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_9 : std_logic_vector (48 to 48);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_7 : std_logic_vector (50 to 50);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_47 : std_logic_vector (10 to 10);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_8 : std_logic_vector (49 to 49);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_44 : std_logic_vector (13 to 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_41 : std_logic_vector (16 to 16);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SALSBS : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_1_0 : std_logic_vector (4 to 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_49_1_0 : std_logic_vector (258 to 258);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M : std_logic_vector (21 downto 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN20_XZXBUS : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2 : std_logic_vector (54 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M14_0X : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M14_0X_0 : std_logic_vector (3 to 3);
  signal GRLFPC2_0_FPO_FRAC : std_logic_vector (54 downto 3);
  signal GRLFPC2_0_COMB_V_I_RES_1 : std_logic_vector (63 downto 29);
  signal GRLFPC2_0_COMB_WRDATA_4 : std_logic_vector (62 downto 0);
  signal GRLFPC2_0_R_I_PC : std_logic_vector (31 downto 2);
  signal GRLFPC2_0_COMB_V_E_STDATA_1 : std_logic_vector (31 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0 : std_logic_vector (56 downto 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_121_0 : std_logic_vector (48 to 48);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT : std_logic_vector (3 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1 : std_logic_vector (56 downto 0);
  signal GRLFPC2_0_COMB_V_I_RES_3 : std_logic_vector (35 downto 32);
  signal GRLFPC2_0_COMB_RS1_1 : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_49_1_2 : std_logic_vector (258 to 258);
  signal GRLFPC2_0_COMB_V_STATE_7 : std_logic_vector (1 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT0 : std_logic_vector (7 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_TZ : std_logic_vector (375 to 375);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_TZ : std_logic_vector (375 to 375);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_129_1 : std_logic_vector (40 to 40);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_130_1 : std_logic_vector (39 to 39);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_149_1 : std_logic_vector (20 to 20);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_135_1 : std_logic_vector (34 to 34);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_150_1 : std_logic_vector (19 to 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_151_1 : std_logic_vector (18 to 18);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_140_1 : std_logic_vector (29 to 29);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_137_1 : std_logic_vector (32 to 32);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_101 : std_logic_vector (12 to 12);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_95 : std_logic_vector (18 to 18);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_111 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_109 : std_logic_vector (4 to 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_108 : std_logic_vector (5 to 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_94 : std_logic_vector (19 to 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_87 : std_logic_vector (26 to 26);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_113 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_64 : std_logic_vector (49 to 49);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_83 : std_logic_vector (30 to 30);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_81 : std_logic_vector (32 to 32);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_80 : std_logic_vector (33 to 33);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_73 : std_logic_vector (40 to 40);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_74 : std_logic_vector (39 to 39);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_85 : std_logic_vector (28 to 28);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_86 : std_logic_vector (27 to 27);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_90 : std_logic_vector (23 to 23);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_106 : std_logic_vector (7 to 7);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_84 : std_logic_vector (29 to 29);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_69 : std_logic_vector (44 to 44);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_98 : std_logic_vector (15 to 15);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_70 : std_logic_vector (43 to 43);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_68 : std_logic_vector (45 to 45);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_67 : std_logic_vector (46 to 46);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_105 : std_logic_vector (8 to 8);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_107 : std_logic_vector (6 to 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_103 : std_logic_vector (10 to 10);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SBLSBS : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SBLSBS_1 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_100 : std_logic_vector (13 to 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_102 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_99 : std_logic_vector (14 to 14);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_97 : std_logic_vector (16 to 16);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_104 : std_logic_vector (9 to 9);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_168_1 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_154_1 : std_logic_vector (15 to 15);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_75 : std_logic_vector (38 to 38);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_76 : std_logic_vector (37 to 37);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_78 : std_logic_vector (35 to 35);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_89 : std_logic_vector (24 to 24);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_88 : std_logic_vector (25 to 25);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_65 : std_logic_vector (48 to 48);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_66 : std_logic_vector (47 to 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE : std_logic_vector (46 downto 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_0 : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_62 : std_logic_vector (51 to 51);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_2_I : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_63 : std_logic_vector (50 to 50);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_0 : std_logic_vector (9 to 9);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_58_1 : std_logic_vector (56 to 56);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_120_1 : std_logic_vector (49 to 49);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0 : std_logic_vector (47 downto 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_1 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_4 : std_logic_vector (3 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL : std_logic_vector (3 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1 : std_logic_vector (7 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_147 : std_logic_vector (22 to 22);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_129 : std_logic_vector (40 to 40);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_130 : std_logic_vector (39 to 39);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_149 : std_logic_vector (20 to 20);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_135 : std_logic_vector (34 to 34);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_150 : std_logic_vector (19 to 19);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_151 : std_logic_vector (18 to 18);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_132 : std_logic_vector (37 to 37);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_164 : std_logic_vector (5 to 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_128 : std_logic_vector (41 to 41);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_140 : std_logic_vector (29 to 29);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_137 : std_logic_vector (32 to 32);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_136 : std_logic_vector (33 to 33);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_145 : std_logic_vector (24 to 24);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_159 : std_logic_vector (10 to 10);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_153 : std_logic_vector (16 to 16);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_167 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_166 : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_165 : std_logic_vector (4 to 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_152 : std_logic_vector (17 to 17);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SCLSBS : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_122 : std_logic_vector (47 to 47);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_139 : std_logic_vector (30 to 30);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_138 : std_logic_vector (31 to 31);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_131 : std_logic_vector (38 to 38);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_143 : std_logic_vector (26 to 26);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_144 : std_logic_vector (25 to 25);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_148 : std_logic_vector (21 to 21);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_156 : std_logic_vector (13 to 13);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_141 : std_logic_vector (28 to 28);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_142 : std_logic_vector (27 to 27);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_155 : std_logic_vector (14 to 14);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_126 : std_logic_vector (43 to 43);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_125 : std_logic_vector (44 to 44);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_127 : std_logic_vector (42 to 42);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_163 : std_logic_vector (6 to 6);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_161 : std_logic_vector (8 to 8);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_168 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_158 : std_logic_vector (11 to 11);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_157 : std_logic_vector (12 to 12);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_160 : std_logic_vector (9 to 9);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_162 : std_logic_vector (7 to 7);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_154 : std_logic_vector (15 to 15);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_133 : std_logic_vector (36 to 36);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_134 : std_logic_vector (35 to 35);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_146 : std_logic_vector (23 to 23);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_1 : std_logic_vector (57 downto 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_123 : std_logic_vector (46 to 46);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_124 : std_logic_vector (45 to 45);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_121 : std_logic_vector (48 to 48);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SCLSBS_1 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14_M_1 : std_logic_vector (171 to 171);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8 : std_logic_vector (57 downto 8);
  signal GRLFPC2_0_R_I_CC : std_logic_vector (1 downto 0);
  signal GRLFPC2_0_COMB_V_FSR_FCC_1_M1 : std_logic_vector (1 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_114_1 : std_logic_vector (56 to 56);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_117 : std_logic_vector (52 to 52);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_3 : std_logic_vector (57 to 57);
  signal GRLFPC2_0_R_A_RF2REN : std_logic_vector (2 downto 1);
  signal GRLFPC2_0_R_A_RF1REN : std_logic_vector (2 downto 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4 : std_logic_vector (57 downto 4);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_2 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2 : std_logic_vector (1 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_I : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8 : std_logic_vector (9 downto 8);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2 : std_logic_vector (56 downto 2);
  signal GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_0 : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_49_1 : std_logic_vector (258 to 258);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8 : std_logic_vector (55 downto 0);
  signal GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_1 : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_5 : std_logic_vector (57 to 57);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_3 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_M : std_logic_vector (21 downto 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_1 : std_logic_vector (57 to 57);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M : std_logic_vector (53 to 53);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M_0 : std_logic_vector (56 downto 8);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH : std_logic_vector (257 downto 58);
  signal GRLFPC2_0_COMB_V_FSR_RD_1 : std_logic_vector (1 downto 0);
  signal GRLFPC2_0_COMB_V_FSR_TEM_1 : std_logic_vector (4 downto 0);
  signal GRLFPC2_0_COMB_V_STATE_1 : std_logic_vector (1 downto 0);
  signal GRLFPC2_0_COMB_V_FSR_FCC_1 : std_logic_vector (1 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_3_I : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23_I_I : std_logic_vector (60 to 60);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_49 : std_logic_vector (258 to 258);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_1_1 : std_logic_vector (57 to 57);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_0_1 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_R_X_RDD_0_0_TMP_D_ARRAY_0 : std_logic_vector (0 to 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_0X : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_0_RN_0 : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS_0_0_0_1 : std_logic_vector (5 to 5);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_1_1 : std_logic_vector (57 to 57);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_M_0_1 : std_logic_vector (7 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M_0_1 : std_logic_vector (44 downto 8);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_0_1 : std_logic_vector (176 to 176);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_2_1_1_0 : std_logic_vector (1 to 1);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_RN_0 : std_logic_vector (2 to 2);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_SN : std_logic_vector (2 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_RN_1 : std_logic_vector (1 downto 0);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_1_0 : std_logic_vector (3 to 3);
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN4_TEMP_2_0_RN_1 : std_logic_vector (0 to 0);
  signal CPO_EXC_INT_2 : std_logic ;
  signal CPO_CC_0_INT_3 : std_logic ;
  signal CPO_CC_1_INT_4 : std_logic ;
  signal RFI2_RD1ADDR_0_INT_5_INT_17 : std_logic ;
  signal RFI2_RD1ADDR_1_INT_6_INT_18 : std_logic ;
  signal RFI2_RD1ADDR_2_INT_7_INT_19 : std_logic ;
  signal RFI2_RD1ADDR_3_INT_8_INT_20 : std_logic ;
  signal RFI2_RD2ADDR_0_INT_9_INT_21 : std_logic ;
  signal RFI2_RD2ADDR_1_INT_10_INT_22 : std_logic ;
  signal RFI2_RD2ADDR_2_INT_11_INT_23 : std_logic ;
  signal RFI2_RD2ADDR_3_INT_12_INT_24 : std_logic ;
  signal RFI2_WRADDR_0_INT_13_INT_25 : std_logic ;
  signal RFI2_WRADDR_1_INT_14_INT_26 : std_logic ;
  signal RFI2_WRADDR_2_INT_15_INT_27 : std_logic ;
  signal RFI2_WRADDR_3_INT_16_INT_28 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1997_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SCTRL_NEW_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1728_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1741_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_760 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_752 : std_logic ;
  signal GRLFPC2_0_N_774_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1723_I : std_logic ;
  signal GRLFPC2_0_FPI_START : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN2_NOTDECODEDUNIMP_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_UN72_PCTRL_NEW_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1519_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTRESETORUNIMP_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_UN61_PCTRL_NEW_I : std_logic ;
  signal NN_1 : std_logic ;
  signal NN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_0_AND : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_1_AND : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_2_AND : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_3_AND : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_4_AND : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_5_AND : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_6_AND : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_7_AND : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT : std_logic ;
  signal GRLFPC2_0_R_I_V : std_logic ;
  signal GRLFPC2_0_COMB_V_I_V_1 : std_logic ;
  signal RST_I : std_logic ;
  signal GRLFPC2_0_V_I_V_3_SQMUXA_I : std_logic ;
  signal GRLFPC2_0_R_MK_BUSY : std_logic ;
  signal GRLFPC2_0_COMB_V_MK_BUSY_2 : std_logic ;
  signal GRLFPC2_0_R_MK_BUSY2 : std_logic ;
  signal GRLFPC2_0_COMB_V_MK_BUSY2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1990_I : std_logic ;
  signal GRLFPC2_0_COMB_UN2_HOLDN : std_logic ;
  signal GRLFPC2_0_N_762_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1996_I : std_logic ;
  signal GRLFPC2_0_R_MK_HOLDN1 : std_logic ;
  signal GRLFPC2_0_R_MK_RST2_I : std_logic ;
  signal N_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_8 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_8 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_9 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_9 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_10 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_10 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_11 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_11 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_12 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_0 : std_logic ;
  signal N_2456 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_1 : std_logic ;
  signal N_2457 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_2 : std_logic ;
  signal N_2458 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_3 : std_logic ;
  signal N_2459 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_4 : std_logic ;
  signal N_2460 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_5 : std_logic ;
  signal N_2461 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_6 : std_logic ;
  signal N_2462 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_7 : std_logic ;
  signal N_2463 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_8 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_8 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_9 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_9 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_998 : std_logic ;
  signal N_2483 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_10 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_10 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_999 : std_logic ;
  signal N_2490 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_11 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_11 : std_logic ;
  signal N_2476 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_12 : std_logic ;
  signal N_2477 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_8 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_8 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_9 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_9 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_10 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_10 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_11 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_11 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_12 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_12 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_13 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_13 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_14 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_14 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_15 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_15 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_16 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_16 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_17 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_17 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_18 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_18 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_19 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_19 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_20 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_20 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_21 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_21 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_22 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_22 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_23 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_23 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_24 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_24 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_25 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_25 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_26 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_26 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_27 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_27 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_28 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_28 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_29 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_29 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_30 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_30 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_31 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_31 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2 : std_logic ;
  signal N_2564 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_32 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_32 : std_logic ;
  signal N_2568 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_33 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_33 : std_logic ;
  signal N_2572 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_34 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_34 : std_logic ;
  signal N_2576 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_35 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_35 : std_logic ;
  signal N_2580 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_36 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_36 : std_logic ;
  signal N_2584 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_37 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_37 : std_logic ;
  signal N_2588 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_38 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_38 : std_logic ;
  signal N_2592 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_39 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_39 : std_logic ;
  signal N_2596 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_40 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_40 : std_logic ;
  signal N_2600 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_41 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_41 : std_logic ;
  signal N_2604 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_42 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_42 : std_logic ;
  signal N_2608 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_43 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_43 : std_logic ;
  signal N_2612 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_44 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_44 : std_logic ;
  signal N_2616 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_45 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_45 : std_logic ;
  signal N_2620 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_46 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_46 : std_logic ;
  signal N_2624 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_47 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_47 : std_logic ;
  signal N_2628 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_48 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_48 : std_logic ;
  signal N_2632 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_49 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_49 : std_logic ;
  signal N_2636 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_50 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_50 : std_logic ;
  signal N_2640 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_51 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_51 : std_logic ;
  signal N_2644 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_52 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_52 : std_logic ;
  signal N_2648 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_53 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_53 : std_logic ;
  signal N_2652 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_54 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_54 : std_logic ;
  signal N_20281 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_55 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_55 : std_logic ;
  signal N_2656 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_56 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_56 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_57 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_8 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_8 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_9 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_9 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_10 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_10 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_11 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_11 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_12 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_12 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_13 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_13 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_14 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_14 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_15 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_15 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_16 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_16 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_17 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_17 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_18 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_18 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_19 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_19 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_20 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_20 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_21 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_21 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_22 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_22 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_23 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_23 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_24 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_24 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_25 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_25 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_26 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_26 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_27 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_27 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_28 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_28 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_29 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_29 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_30 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_30 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_31 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_31 : std_logic ;
  signal N_2724 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_32 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_32 : std_logic ;
  signal N_2731 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_33 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_33 : std_logic ;
  signal N_2738 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_34 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_34 : std_logic ;
  signal N_2745 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_35 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_35 : std_logic ;
  signal N_2752 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_36 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_36 : std_logic ;
  signal N_2759 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_37 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_37 : std_logic ;
  signal N_2766 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_38 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_38 : std_logic ;
  signal N_2773 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_39 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_39 : std_logic ;
  signal N_2780 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_40 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_40 : std_logic ;
  signal N_2787 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_41 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_41 : std_logic ;
  signal N_2794 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_42 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_42 : std_logic ;
  signal N_2801 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_43 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_43 : std_logic ;
  signal N_2808 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_44 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_44 : std_logic ;
  signal N_2815 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_45 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_45 : std_logic ;
  signal N_2822 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_46 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_46 : std_logic ;
  signal N_2829 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_47 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_47 : std_logic ;
  signal N_2836 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_48 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_48 : std_logic ;
  signal N_2843 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_49 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_49 : std_logic ;
  signal N_2850 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_50 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_50 : std_logic ;
  signal N_2857 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_51 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_51 : std_logic ;
  signal N_2864 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_52 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_52 : std_logic ;
  signal N_2871 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_53 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_53 : std_logic ;
  signal N_2878 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_54 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_54 : std_logic ;
  signal N_20279 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_55 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_55 : std_logic ;
  signal N_2885 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_56 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_56 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_57 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2032_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN20_U_RDN_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1749_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1748_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_115_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELECTDIVMULT_UN86_DIVMULTV : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2297 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2298 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_814 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_815 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_813 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_812 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_811 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_810 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_113_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_112_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_111_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_110_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_109_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_108_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_107_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_106_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_105_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_104_I : std_logic ;
  signal N_8694_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2342 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_102_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_101_I : std_logic ;
  signal N_8699_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2207 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_99_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_98_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_97_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_96_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_95_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_94_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_93_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_92_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_91_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_90_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_89_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_88_I : std_logic ;
  signal N_8692_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2338 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_86_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_85_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_84_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_83_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_82_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_81_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_80_I : std_logic ;
  signal N_8693_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2323 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_78_I : std_logic ;
  signal N_8688_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2328 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_76_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_75_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_74_I : std_logic ;
  signal N_8689_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2334 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_72_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_71_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_70_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_69_I : std_logic ;
  signal N_8700_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2302 : std_logic ;
  signal N_8690_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2305 : std_logic ;
  signal N_8701_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2309 : std_logic ;
  signal N_8691_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2312 : std_logic ;
  signal N_8702_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2316 : std_logic ;
  signal N_8687_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2319 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_62_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_61_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_60_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_59_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_58_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_57_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_0 : std_logic ;
  signal N_8703_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2299 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_55_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_54_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_53_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_52_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_51_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_50_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_49_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_48_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_47_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_46_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_45_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_44_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_43_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_42_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_41_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_40_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_39_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_38_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_37_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_36_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_35_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_34_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_33_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_32_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_31_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_30_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_29_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_28_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_27_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_26_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_25_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_24_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_23_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_22_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_21_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_20_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_19_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_18_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_17_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_16_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_15_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_14_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_13_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_12_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_11_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_10_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_9_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_8_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_7_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_6_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_5_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_4_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_3_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_2_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_1_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_0_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_I : std_logic ;
  signal GRLFPC2_0_R_MK_LDOP : std_logic ;
  signal GRLFPC2_0_R_MK_LDOPC : std_logic ;
  signal GRLFPC2_0_R_MK_RST : std_logic ;
  signal GRLFPC2_0_R_MK_RSTC : std_logic ;
  signal HOLDN_I : std_logic ;
  signal GRLFPC2_0_COMB_RS2_1_SN_N_2 : std_logic ;
  signal N_6758 : std_logic ;
  signal N_6759 : std_logic ;
  signal N_6760 : std_logic ;
  signal N_6761 : std_logic ;
  signal N_6762 : std_logic ;
  signal N_6763 : std_logic ;
  signal N_6764 : std_logic ;
  signal N_6765 : std_logic ;
  signal N_6766 : std_logic ;
  signal N_6767 : std_logic ;
  signal N_6768 : std_logic ;
  signal N_6769 : std_logic ;
  signal N_6770 : std_logic ;
  signal N_6771 : std_logic ;
  signal N_6772 : std_logic ;
  signal N_6773 : std_logic ;
  signal N_6774 : std_logic ;
  signal N_6775 : std_logic ;
  signal N_6776 : std_logic ;
  signal N_6777 : std_logic ;
  signal N_6778 : std_logic ;
  signal N_6779 : std_logic ;
  signal N_6780 : std_logic ;
  signal N_6781 : std_logic ;
  signal N_6782 : std_logic ;
  signal N_6783 : std_logic ;
  signal N_6784 : std_logic ;
  signal N_6785 : std_logic ;
  signal N_6786 : std_logic ;
  signal N_6787 : std_logic ;
  signal N_6788 : std_logic ;
  signal N_6789 : std_logic ;
  signal N_6790 : std_logic ;
  signal N_6791 : std_logic ;
  signal N_6792 : std_logic ;
  signal N_6793 : std_logic ;
  signal N_6794 : std_logic ;
  signal N_6795 : std_logic ;
  signal N_6796 : std_logic ;
  signal N_6797 : std_logic ;
  signal N_6798 : std_logic ;
  signal N_6799 : std_logic ;
  signal N_6800 : std_logic ;
  signal N_6801 : std_logic ;
  signal N_6802 : std_logic ;
  signal N_6803 : std_logic ;
  signal N_6804 : std_logic ;
  signal N_6805 : std_logic ;
  signal N_6806 : std_logic ;
  signal N_6807 : std_logic ;
  signal N_6808 : std_logic ;
  signal N_6809 : std_logic ;
  signal N_6810 : std_logic ;
  signal N_6811 : std_logic ;
  signal N_6812 : std_logic ;
  signal N_6813 : std_logic ;
  signal N_6814 : std_logic ;
  signal N_6815 : std_logic ;
  signal N_6816 : std_logic ;
  signal N_6817 : std_logic ;
  signal N_6818 : std_logic ;
  signal N_6819 : std_logic ;
  signal N_6820 : std_logic ;
  signal N_6829_A : std_logic ;
  signal N_6830_A : std_logic ;
  signal N_6831_A : std_logic ;
  signal N_6832_A : std_logic ;
  signal N_6833_A : std_logic ;
  signal N_6834_A : std_logic ;
  signal N_6835_A : std_logic ;
  signal N_6836_A : std_logic ;
  signal N_6837_A : std_logic ;
  signal N_6838_A : std_logic ;
  signal N_6839_A : std_logic ;
  signal N_6840_A : std_logic ;
  signal N_6841_A : std_logic ;
  signal N_6842_A : std_logic ;
  signal N_6843_A : std_logic ;
  signal N_6844_A : std_logic ;
  signal N_6845_A : std_logic ;
  signal N_6846_A : std_logic ;
  signal N_6847_A : std_logic ;
  signal N_6848_A : std_logic ;
  signal N_6849_A : std_logic ;
  signal N_6850_A : std_logic ;
  signal N_6851_A : std_logic ;
  signal N_6852_A : std_logic ;
  signal N_6853_A : std_logic ;
  signal N_6854_A : std_logic ;
  signal N_6855_A : std_logic ;
  signal N_6856_A : std_logic ;
  signal N_6857_A : std_logic ;
  signal N_6858_A : std_logic ;
  signal N_6859_A : std_logic ;
  signal N_6860_A : std_logic ;
  signal N_6861_A : std_logic ;
  signal N_6862_A : std_logic ;
  signal N_6863_A : std_logic ;
  signal N_6864_A : std_logic ;
  signal N_6865_A : std_logic ;
  signal N_6866_A : std_logic ;
  signal N_6867_A : std_logic ;
  signal N_6868_A : std_logic ;
  signal N_6869_A : std_logic ;
  signal N_6870_A : std_logic ;
  signal N_6871_A : std_logic ;
  signal N_6872_A : std_logic ;
  signal N_6873_A : std_logic ;
  signal N_6874_A : std_logic ;
  signal N_6875_A : std_logic ;
  signal N_6876_A : std_logic ;
  signal N_6877_A : std_logic ;
  signal N_6878_A : std_logic ;
  signal N_6879_A : std_logic ;
  signal N_6880_A : std_logic ;
  signal N_6881_A : std_logic ;
  signal N_6882_A : std_logic ;
  signal N_6883_A : std_logic ;
  signal N_6884_A : std_logic ;
  signal N_6885_A : std_logic ;
  signal N_6886_A : std_logic ;
  signal N_6887_A : std_logic ;
  signal N_6888_A : std_logic ;
  signal N_6889_A : std_logic ;
  signal N_6890_A : std_logic ;
  signal N_6891_A : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SM3_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2030 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_ROMXZSL2FROMC : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_7_AND1 : std_logic ;
  signal GRLFPC2_0_R_MK_HOLDN2 : std_logic ;
  signal GRLFPC2_0_R_MK_RST2 : std_logic ;
  signal GRLFPC2_0_N_782 : std_logic ;
  signal GRLFPC2_0_SEQERR_1_SQMUXA_1_SN : std_logic ;
  signal GRLFPC2_0_MOV_0_SQMUXA_2 : std_logic ;
  signal GRLFPC2_0_MOV_2_SQMUXA_2 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_MOV6_2 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_AFQ12 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_AFQ13 : std_logic ;
  signal GRLFPC2_0_COMB_V_E_STDATA2 : std_logic ;
  signal GRLFPC2_0_R_M_FPOP : std_logic ;
  signal GRLFPC2_0_COMB_UN22_CCV : std_logic ;
  signal GRLFPC2_0_R_X_FPOP : std_logic ;
  signal GRLFPC2_0_COMB_UN14_CCV : std_logic ;
  signal GRLFPC2_0_R_E_FPOP : std_logic ;
  signal GRLFPC2_0_ANNULRES_0_SQMUXA_3_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_AREGXORBREG : std_logic ;
  signal GRLFPC2_0_R_X_AFSR : std_logic ;
  signal GRLFPC2_0_R_X_LD : std_logic ;
  signal GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA : std_logic ;
  signal GRLFPC2_0_COMB_WREN22 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2031 : std_logic ;
  signal GRLFPC2_0_N_703_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SM6_I : std_logic ;
  signal GRLFPC2_0_MOV_2_SQMUXA_1_0 : std_logic ;
  signal GRLFPC2_0_MOV_0_SQMUXA_3 : std_logic ;
  signal GRLFPC2_0_COMB_UN1_FPCI_1_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2281_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_ENTRYSHFT_S_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN19_FEEDBACK_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SM0_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_16_REP1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN23_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV_4_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN5_NOTSHIFTCOUNT1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_2_SN_M1_E_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_992 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1000 : std_logic ;
  signal GRLFPC2_0_N_311 : std_logic ;
  signal GRLFPC2_0_N_312 : std_logic ;
  signal GRLFPC2_0_N_313 : std_logic ;
  signal GRLFPC2_0_N_314 : std_logic ;
  signal GRLFPC2_0_N_316 : std_logic ;
  signal GRLFPC2_0_N_317 : std_logic ;
  signal GRLFPC2_0_N_318 : std_logic ;
  signal GRLFPC2_0_N_319 : std_logic ;
  signal GRLFPC2_0_N_320 : std_logic ;
  signal GRLFPC2_0_N_321 : std_logic ;
  signal GRLFPC2_0_N_322 : std_logic ;
  signal GRLFPC2_0_N_333 : std_logic ;
  signal GRLFPC2_0_N_334 : std_logic ;
  signal GRLFPC2_0_N_335 : std_logic ;
  signal GRLFPC2_0_N_336 : std_logic ;
  signal GRLFPC2_0_N_338 : std_logic ;
  signal GRLFPC2_0_N_341 : std_logic ;
  signal GRLFPC2_0_N_342 : std_logic ;
  signal GRLFPC2_0_N_325 : std_logic ;
  signal GRLFPC2_0_N_315 : std_logic ;
  signal GRLFPC2_0_N_337 : std_logic ;
  signal GRLFPC2_0_N_327 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELINITREMBIT : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2017 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2016 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_COMPUTECONST_UN49_RESVEC : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_NOTAM2_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN19_FEEDBACK : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_3_SN_I3_I_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2003 : std_logic ;
  signal GRLFPC2_0_R_I_EXEC : std_logic ;
  signal GRLFPC2_0_COMB_UN1_R_I_V : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_AFQ4_1 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_AFQ7_1 : std_logic ;
  signal GRLFPC2_0_MOV_7_SQMUXA_3 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_MOV5_1 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_1_0 : std_logic ;
  signal GRLFPC2_0_ANNULFPU_0_SQMUXA_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_854 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTXZYFROMD_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_2_0 : std_logic ;
  signal GRLFPC2_0_R_MK_LDOPC_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN9_S_11_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_53_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN11_NOTBINFNAN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN11_NOTAINFNAN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN5_NOTBZERODENORM_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN5_NOTAZERODENORM_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN5_XZYBUSLSBS : std_logic ;
  signal GRLFPC2_0_N_781 : std_logic ;
  signal GRLFPC2_0_R_A_LD : std_logic ;
  signal GRLFPC2_0_R_E_LD : std_logic ;
  signal GRLFPC2_0_R_M_LD : std_logic ;
  signal GRLFPC2_0_N_776 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_RS2D5_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN18_FEEDBACK : std_logic ;
  signal GRLFPC2_0_R_A_RS1D : std_logic ;
  signal GRLFPC2_0_R_A_ST : std_logic ;
  signal GRLFPC2_0_COMB_UN1_FPCI_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_6_AND_1 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_AFQ8_0 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_UN1_WREN210_1_0_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_S_CMP_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN14_S_MOV_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTAINFNAN_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTAINFNAN_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTBINFNAN_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTBINFNAN_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_I_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_I_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV_6_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN17_SRTOSTICKY_3 : std_logic ;
  signal GRLFPC2_0_R_MK_LDOPC_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_UN525_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_UN354_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_UN183_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_UN12_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_UN363_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_UN534_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_UN573_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_UN402_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_UN231_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_UN60_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_UN636_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_UN465_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_UN294_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_UN123_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2008 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_UN540_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_UN369_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_UN198_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_UN639_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_UN468_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_UN297_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_UN126_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_UN129_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_UN300_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_UN471_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_UN642_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_UN168_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_UN633_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_19_TRFWWBASICCELL_UN624_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_UN462_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_UN291_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_UN120_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_19_TRFWWBASICCELL_UN111_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_UN597_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_UN426_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_UN255_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_UN84_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_UN510_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_UN339_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_UN651_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_UN480_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_UN309_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_UN138_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_UN648_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_UN477_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_UN306_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_UN135_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_UN3_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_UN6_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_UN9_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_UN15_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_UN18_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_UN30_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_UN33_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_UN36_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_UN39_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_UN42_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_UN45_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_UN48_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_UN51_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_UN54_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_UN57_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_UN63_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_UN66_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_UN69_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_UN72_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_UN75_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_UN78_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_UN81_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_UN87_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_UN90_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_UN93_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_UN96_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_UN99_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_UN102_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_UN105_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_UN108_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_18_TRFWWBASICCELL_UN114_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_UN117_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_UN132_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_UN141_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_UN144_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_UN147_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_UN150_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_UN153_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_UN156_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_UN159_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_UN162_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_UN165_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_UN171_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_UN174_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_UN177_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_UN180_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_UN186_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_UN201_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_UN204_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_UN207_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_UN210_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_UN216_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_UN219_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_UN222_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_UN225_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_UN228_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_UN234_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_UN237_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_UN240_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_UN243_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_UN246_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_UN252_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_UN258_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_UN261_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_UN264_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_UN267_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_UN270_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_UN273_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_UN276_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_UN288_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_UN303_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_UN312_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_UN315_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_UN318_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_UN321_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_UN324_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_UN327_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_UN330_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_UN333_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_UN336_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_UN342_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_UN345_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_UN348_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_UN351_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_UN357_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_UN360_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_UN366_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_UN372_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_UN375_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_UN378_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_UN381_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_UN384_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_UN387_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_UN390_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_UN393_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_UN396_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_UN399_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_UN405_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_UN408_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_UN411_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_UN414_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_UN417_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_UN420_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_UN423_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_UN429_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_UN432_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_UN435_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_UN438_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_UN441_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_UN444_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_UN447_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_UN450_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_UN459_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_UN474_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_UN483_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_UN486_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_UN489_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_UN492_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_UN495_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_UN498_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_UN501_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_UN504_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_UN507_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_UN513_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_UN516_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_UN519_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_UN522_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_UN528_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_UN531_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_UN537_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_UN543_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_UN546_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_UN549_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_UN552_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_UN555_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_UN558_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_UN561_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_UN570_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_UN576_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_UN579_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_UN582_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_UN585_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_UN588_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_UN591_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_UN594_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_UN600_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_UN603_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_UN606_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_UN609_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_UN612_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_UN615_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_UN618_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_UN621_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_18_TRFWWBASICCELL_UN627_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_UN630_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_UN645_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_UN654_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_UN657_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_UN660_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_UN663_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_UN666_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_UN669_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_UN672_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_UN675_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_UN678_TEMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SS6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_846 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1017 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_42_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_44_0 : std_logic ;
  signal GRLFPC2_0_R_X_AFQ : std_logic ;
  signal GRLFPC2_0_R_X_SEQERR : std_logic ;
  signal GRLFPC2_0_V_STATE_1_SQMUXA_1 : std_logic ;
  signal GRLFPC2_0_V_FSR_FTT_1_SQMUXA_2_2 : std_logic ;
  signal GRLFPC2_0_WREN2_1_SQMUXA_1 : std_logic ;
  signal GRLFPC2_0_V_I_EXEC_0_SQMUXA : std_logic ;
  signal GRLFPC2_0_WRADDR_0_SQMUXA_1 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_UN3_OP : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_AFQ3 : std_logic ;
  signal GRLFPC2_0_N_772 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CONDMUXMULXFF_UN4_NOTSQRTLFTCC : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_AFQ7 : std_logic ;
  signal GRLFPC2_0_V_FSR_AEXC_1_SQMUXA_SN : std_logic ;
  signal GRLFPC2_0_R_A_RS2D : std_logic ;
  signal GRLFPC2_0_N_771 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN46_XZYBUSLSBS : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN3_INEXACT : std_logic ;
  signal N_12084 : std_logic ;
  signal GRLFPC2_0_R_FSR_NONSTD : std_logic ;
  signal N_12086 : std_logic ;
  signal N_12087 : std_logic ;
  signal GRLFPC2_0_R_A_FPOP : std_logic ;
  signal GRLFPC2_0_ANNULRES_0_SQMUXA_3_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN1_MIFROMINST_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0 : std_logic ;
  signal GRLFPC2_0_R_A_MOV : std_logic ;
  signal GRLFPC2_0_N_691 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_S_CMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1991 : std_logic ;
  signal GRLFPC2_0_N_777 : std_logic ;
  signal GRLFPC2_0_MOV_2_SQMUXA_1_1 : std_logic ;
  signal GRLFPC2_0_COMB_UN8_CCV_1 : std_logic ;
  signal GRLFPC2_0_COMB_LOCK_1_1_0 : std_logic ;
  signal GRLFPC2_0_COMB_ANNULFPU_1_U_0 : std_logic ;
  signal GRLFPC2_0_COMB_UN1_MEXC_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN4_S_SQRT_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_845 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_847 : std_logic ;
  signal N_12088 : std_logic ;
  signal N_12089 : std_logic ;
  signal N_12090 : std_logic ;
  signal N_12091 : std_logic ;
  signal N_12092 : std_logic ;
  signal N_12093 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1019 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1020 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1021 : std_logic ;
  signal GRLFPC2_0_COMB_ISFPOP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_844 : std_logic ;
  signal GRLFPC2_0_N_206 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_16_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_23_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_19_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN39_XZYBUSLSBS : std_logic ;
  signal GRLFPC2_0_N_716 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN1_U_SNNOTDB : std_logic ;
  signal GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1 : std_logic ;
  signal GRLFPC2_0_V_STATE_1_SQMUXA : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN12_U_SNNOTDB_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2000 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_18_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_18_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_TEMP2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_19_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_TEMP2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_19_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_TEMP2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_TEMP2_1 : std_logic ;
  signal N_5258 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_MOV5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_12_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_11_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_10_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN14_S_MOV : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2002 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTBINFNAN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTAINFNAN : std_logic ;
  signal GRLFPC2_0_MOV_7_SQMUXA : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_RS2D5_3 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_RS2D5 : std_logic ;
  signal GRLFPC2_0_COMB_UN6_IUEXEC : std_logic ;
  signal GRLFPC2_0_WREN2_2_SQMUXA : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_MOV6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2023 : std_logic ;
  signal GRLFPC2_0_MOV_5_SQMUXA_2 : std_logic ;
  signal GRLFPC2_0_MOV_0_SQMUXA_2_0 : std_logic ;
  signal GRLFPC2_0_V_STATE_1_SQMUXA_3_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_ENTRYPOINT_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN9_NOTPROP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO : std_logic ;
  signal GRLFPC2_0_COMB_V_FSR_NONSTD_1_M1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SS12 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_104 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_114 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_115 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_116 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_117 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_118 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_119 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_120 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_121 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_122 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_123 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_125 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_126 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_127 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_128 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_129 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_132 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_133 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_134 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_135 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_137 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_138 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_139 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_140 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_141 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_142 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_143 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_144 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_145 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_146 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_147 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_148 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_149 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_150 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_154 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_156 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_157 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_158 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_159 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_161 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_162 : std_logic ;
  signal N_12094 : std_logic ;
  signal N_12095 : std_logic ;
  signal N_12096 : std_logic ;
  signal N_12097 : std_logic ;
  signal N_12098 : std_logic ;
  signal N_12099 : std_logic ;
  signal N_12100 : std_logic ;
  signal N_12101 : std_logic ;
  signal N_12102 : std_logic ;
  signal N_12103 : std_logic ;
  signal N_12104 : std_logic ;
  signal N_12105 : std_logic ;
  signal GRLFPC2_0_N_126 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_155 : std_logic ;
  signal N_12106 : std_logic ;
  signal N_12107 : std_logic ;
  signal N_12108 : std_logic ;
  signal N_12109 : std_logic ;
  signal GRLFPC2_0_N_634 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_163 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_153 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_113 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_124 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_131 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_130 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_136 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_151 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_160 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_152 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN57_SHDVAR : std_logic ;
  signal GRLFPC2_0_N_755 : std_logic ;
  signal GRLFPC2_0_N_653 : std_logic ;
  signal GRLFPC2_0_RS1V10_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24 : std_logic ;
  signal GRLFPC2_0_RS2_0_SQMUXA : std_logic ;
  signal GRLFPC2_0_COMB_SEQERR_UN13_OP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1990 : std_logic ;
  signal N_12110 : std_logic ;
  signal N_12111 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV_6 : std_logic ;
  signal N_12112 : std_logic ;
  signal N_12113 : std_logic ;
  signal N_12114 : std_logic ;
  signal N_12115 : std_logic ;
  signal N_12116 : std_logic ;
  signal N_12117 : std_logic ;
  signal N_12118 : std_logic ;
  signal N_12119 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_353 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN17_WQSTSETS : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP_1 : std_logic ;
  signal GRLFPC2_0_AFQ_3_SQMUXA : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26 : std_logic ;
  signal GRLFPC2_0_WREN2_1_SQMUXA_1_0 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_UN1_WREN210 : std_logic ;
  signal N_2291_TZ : std_logic ;
  signal GRLFPC2_0_COMB_RSDECODE_RS1V2_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA_M1_E_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_N_635 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_19_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_18_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_19_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_CIN_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_CIN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_18_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_CIN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_CIN : std_logic ;
  signal GRLFPC2_0_R_I_RDD : std_logic ;
  signal GRLFPC2_0_R_X_RDD : std_logic ;
  signal GRLFPC2_0_COMB_RDD_3 : std_logic ;
  signal GRLFPC2_0_N_673 : std_logic ;
  signal GRLFPC2_0_COMB_RS1D_1_M1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4 : std_logic ;
  signal GRLFPC2_0_N_710 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_NE_0 : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_MOV11 : std_logic ;
  signal GRLFPC2_0_MOV_3_SQMUXA_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_OPREXCSHFT_UN3_OPREXC : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN42_CONDITIONAL : std_logic ;
  signal GRLFPC2_0_N_766 : std_logic ;
  signal GRLFPC2_0_UN1_AFQ6_I : std_logic ;
  signal GRLFPC2_0_COMB_SEQERR_UN7_OP_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_110 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_111 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_112 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_377 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_378 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_380 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_381 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_383 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_384 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_763 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_764 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_765 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_766 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_768 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_769 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_770 : std_logic ;
  signal GRLFPC2_0_WRADDR_0_SQMUXA : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_382 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_379 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_767 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN1_S_14 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN1_ENTRYPOINT : std_logic ;
  signal GRLFPC2_0_N_764 : std_logic ;
  signal GRLFPC2_0_MOV_2_SQMUXA : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN24_SHDVAR : std_logic ;
  signal GRLFPC2_0_UN1_AFQ7_I_A2_0 : std_logic ;
  signal GRLFPC2_0_RS1V_1_SQMUXA : std_logic ;
  signal GRLFPC2_0_UN1_WREN210_4_0 : std_logic ;
  signal GRLFPC2_0_COMB_V_I_V6_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_ENTRYPOINT_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1870 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2122_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_8 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_9 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_98_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_61_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_88_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_62_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_74_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_96_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_64_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_100_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_78_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_104_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_66_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_94_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_13_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_114_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_NE_2 : std_logic ;
  signal GRLFPC2_0_N_791 : std_logic ;
  signal N_12120 : std_logic ;
  signal N_12121 : std_logic ;
  signal N_12122 : std_logic ;
  signal N_12123 : std_logic ;
  signal N_12124 : std_logic ;
  signal N_12125 : std_logic ;
  signal N_12126 : std_logic ;
  signal N_12127 : std_logic ;
  signal N_12128 : std_logic ;
  signal N_12129 : std_logic ;
  signal N_12130 : std_logic ;
  signal N_12131 : std_logic ;
  signal N_12132 : std_logic ;
  signal N_12133 : std_logic ;
  signal N_12134 : std_logic ;
  signal N_12135 : std_logic ;
  signal N_12136 : std_logic ;
  signal N_12137 : std_logic ;
  signal N_12138 : std_logic ;
  signal N_12139 : std_logic ;
  signal N_12140 : std_logic ;
  signal N_12141 : std_logic ;
  signal N_12142 : std_logic ;
  signal N_12143 : std_logic ;
  signal N_12144 : std_logic ;
  signal N_12145 : std_logic ;
  signal N_12146 : std_logic ;
  signal N_12147 : std_logic ;
  signal N_12148 : std_logic ;
  signal N_12149 : std_logic ;
  signal N_12150 : std_logic ;
  signal N_12151 : std_logic ;
  signal N_12152 : std_logic ;
  signal N_12153 : std_logic ;
  signal N_12154 : std_logic ;
  signal N_12155 : std_logic ;
  signal N_12156 : std_logic ;
  signal N_12157 : std_logic ;
  signal N_12158 : std_logic ;
  signal N_12159 : std_logic ;
  signal N_12160 : std_logic ;
  signal N_12161 : std_logic ;
  signal N_12162 : std_logic ;
  signal N_12163 : std_logic ;
  signal N_12165 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_225 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_279 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2276 : std_logic ;
  signal N_12166 : std_logic ;
  signal N_12167 : std_logic ;
  signal N_12168 : std_logic ;
  signal N_12169 : std_logic ;
  signal N_12170 : std_logic ;
  signal N_12171 : std_logic ;
  signal N_12172 : std_logic ;
  signal N_12173 : std_logic ;
  signal N_12174 : std_logic ;
  signal N_12175 : std_logic ;
  signal N_12176 : std_logic ;
  signal N_12177 : std_logic ;
  signal N_12178 : std_logic ;
  signal N_12179 : std_logic ;
  signal N_12180 : std_logic ;
  signal N_12181 : std_logic ;
  signal GRLFPC2_0_R_A_AFSR : std_logic ;
  signal N_12182 : std_logic ;
  signal N_12183 : std_logic ;
  signal GRLFPC2_0_R_A_AFQ : std_logic ;
  signal N_12184 : std_logic ;
  signal N_12185 : std_logic ;
  signal N_12186 : std_logic ;
  signal N_12187 : std_logic ;
  signal N_12188 : std_logic ;
  signal N_12189 : std_logic ;
  signal N_12190 : std_logic ;
  signal N_12191 : std_logic ;
  signal N_12192 : std_logic ;
  signal N_12193 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_224 : std_logic ;
  signal N_12194 : std_logic ;
  signal N_12195 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_223 : std_logic ;
  signal N_12196 : std_logic ;
  signal N_12197 : std_logic ;
  signal N_12198 : std_logic ;
  signal N_12199 : std_logic ;
  signal N_12200 : std_logic ;
  signal N_12201 : std_logic ;
  signal N_12202 : std_logic ;
  signal N_12203 : std_logic ;
  signal N_12204 : std_logic ;
  signal N_12205 : std_logic ;
  signal N_12206 : std_logic ;
  signal N_12207 : std_logic ;
  signal N_12208 : std_logic ;
  signal N_12209 : std_logic ;
  signal N_12210 : std_logic ;
  signal N_12211 : std_logic ;
  signal N_12212 : std_logic ;
  signal N_12213 : std_logic ;
  signal N_12214 : std_logic ;
  signal N_12215 : std_logic ;
  signal N_12216 : std_logic ;
  signal N_12217 : std_logic ;
  signal GRLFPC2_0_COMB_V_I_V6 : std_logic ;
  signal GRLFPC2_0_COMB_WREN2_9_IV_0 : std_logic ;
  signal N_12218 : std_logic ;
  signal N_12219 : std_logic ;
  signal N_12220 : std_logic ;
  signal N_12221 : std_logic ;
  signal N_12222 : std_logic ;
  signal N_12223 : std_logic ;
  signal N_12224 : std_logic ;
  signal N_12225 : std_logic ;
  signal N_12226 : std_logic ;
  signal N_12227 : std_logic ;
  signal N_12228 : std_logic ;
  signal N_12229 : std_logic ;
  signal N_12230 : std_logic ;
  signal N_12231 : std_logic ;
  signal N_12232 : std_logic ;
  signal N_12233 : std_logic ;
  signal N_12234 : std_logic ;
  signal N_12235 : std_logic ;
  signal N_12236 : std_logic ;
  signal N_12237 : std_logic ;
  signal N_12238 : std_logic ;
  signal N_12239 : std_logic ;
  signal N_12240 : std_logic ;
  signal N_12241 : std_logic ;
  signal N_12242 : std_logic ;
  signal N_12243 : std_logic ;
  signal N_12244 : std_logic ;
  signal N_12245 : std_logic ;
  signal N_12246 : std_logic ;
  signal N_12247 : std_logic ;
  signal N_12248 : std_logic ;
  signal N_12249 : std_logic ;
  signal N_12250 : std_logic ;
  signal N_12251 : std_logic ;
  signal N_12252 : std_logic ;
  signal N_12253 : std_logic ;
  signal N_12254 : std_logic ;
  signal N_12255 : std_logic ;
  signal N_12256 : std_logic ;
  signal N_12257 : std_logic ;
  signal GRLFPC2_0_UN1_AFQ3_I : std_logic ;
  signal GRLFPC2_0_COMB_RS1D_1_M2 : std_logic ;
  signal GRLFPC2_0_N_674 : std_logic ;
  signal N_12258 : std_logic ;
  signal N_12259 : std_logic ;
  signal N_12260 : std_logic ;
  signal N_12261 : std_logic ;
  signal N_12262 : std_logic ;
  signal N_12263 : std_logic ;
  signal N_8928 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_15 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT : std_logic ;
  signal GRLFPC2_0_N_670 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_NE_4 : std_logic ;
  signal GRLFPC2_0_V_STATE_2_SQMUXA : std_logic ;
  signal GRLFPC2_0_N_789 : std_logic ;
  signal GRLFPC2_0_V_FSR_FTT_1_SQMUXA_2_1 : std_logic ;
  signal GRLFPC2_0_N_736 : std_logic ;
  signal GRLFPC2_0_V_I_EXEC26 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_0 : std_logic ;
  signal N_12264 : std_logic ;
  signal N_12265 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1549 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1550 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1551 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1552 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1546 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1547 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1548 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1542 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1543 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1544 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1545 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1539 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1537 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1571 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1566 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1567 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1561 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1557 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1559 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1560 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1553 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1554 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1555 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1556 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1579 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1580 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1581 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1576 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1577 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1573 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1575 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1569 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1570 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1583 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1585 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTDECODEDUNIMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1533 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1535 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1534 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1541 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1540 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1538 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1565 : std_logic ;
  signal GRLFPC2_0_UN1_AFQ7_I_A2_2 : std_logic ;
  signal GRLFPC2_0_COMB_RDD_1_0_0 : std_logic ;
  signal GRLFPC2_0_COMB_V_A_AFSR_1_0_1 : std_logic ;
  signal GRLFPC2_0_I_162_1 : std_logic ;
  signal GRLFPC2_0_COMB_RS1D_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_71 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1935 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1949 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1948 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1945 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1942 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1940 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1939 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1965 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1964 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1963 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1962 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1960 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1959 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1957 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1956 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1955 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1953 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1952 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1980 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1977 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1983 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1982 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1934 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1958 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1978 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1979 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1981 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1987 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1967 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1966 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1943 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1944 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1950 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1951 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1954 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1936 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1937 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1961 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1973 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1974 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1938 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1941 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1968 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1969 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1970 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1971 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1972 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1984 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1985 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1975 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1976 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1947 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1946 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_278 : std_logic ;
  signal N_12266 : std_logic ;
  signal N_12267 : std_logic ;
  signal N_12268 : std_logic ;
  signal N_12269 : std_logic ;
  signal N_12270 : std_logic ;
  signal N_12271 : std_logic ;
  signal N_12272 : std_logic ;
  signal N_12273 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_363 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_566 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_568 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_569 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_570 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_571 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_573 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_574 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_575 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_576 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_577 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_585 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_586 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_588 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_590 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_596 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_599 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_601 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_603 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_604 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_605 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_607 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_609 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_610 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_615 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_616 : std_logic ;
  signal GRLFPC2_0_N_63 : std_logic ;
  signal GRLFPC2_0_N_65 : std_logic ;
  signal GRLFPC2_0_N_67 : std_logic ;
  signal GRLFPC2_0_N_68 : std_logic ;
  signal GRLFPC2_0_N_69 : std_logic ;
  signal GRLFPC2_0_N_70 : std_logic ;
  signal GRLFPC2_0_N_71 : std_logic ;
  signal GRLFPC2_0_N_72 : std_logic ;
  signal GRLFPC2_0_N_73 : std_logic ;
  signal GRLFPC2_0_N_74 : std_logic ;
  signal GRLFPC2_0_N_75 : std_logic ;
  signal GRLFPC2_0_N_77 : std_logic ;
  signal GRLFPC2_0_N_78 : std_logic ;
  signal GRLFPC2_0_N_81 : std_logic ;
  signal GRLFPC2_0_N_82 : std_logic ;
  signal GRLFPC2_0_N_84 : std_logic ;
  signal GRLFPC2_0_N_85 : std_logic ;
  signal GRLFPC2_0_N_86 : std_logic ;
  signal GRLFPC2_0_N_87 : std_logic ;
  signal GRLFPC2_0_N_88 : std_logic ;
  signal GRLFPC2_0_N_89 : std_logic ;
  signal GRLFPC2_0_N_91 : std_logic ;
  signal GRLFPC2_0_N_92 : std_logic ;
  signal GRLFPC2_0_N_94 : std_logic ;
  signal GRLFPC2_0_N_95 : std_logic ;
  signal GRLFPC2_0_N_97 : std_logic ;
  signal GRLFPC2_0_N_99 : std_logic ;
  signal GRLFPC2_0_N_100 : std_logic ;
  signal GRLFPC2_0_N_101 : std_logic ;
  signal GRLFPC2_0_N_102 : std_logic ;
  signal GRLFPC2_0_N_103 : std_logic ;
  signal GRLFPC2_0_N_104 : std_logic ;
  signal GRLFPC2_0_N_105 : std_logic ;
  signal GRLFPC2_0_N_106 : std_logic ;
  signal GRLFPC2_0_N_107 : std_logic ;
  signal GRLFPC2_0_N_109 : std_logic ;
  signal GRLFPC2_0_N_110 : std_logic ;
  signal GRLFPC2_0_N_113 : std_logic ;
  signal GRLFPC2_0_N_114 : std_logic ;
  signal GRLFPC2_0_N_116 : std_logic ;
  signal GRLFPC2_0_N_117 : std_logic ;
  signal GRLFPC2_0_N_118 : std_logic ;
  signal GRLFPC2_0_N_119 : std_logic ;
  signal GRLFPC2_0_N_120 : std_logic ;
  signal GRLFPC2_0_N_121 : std_logic ;
  signal GRLFPC2_0_N_123 : std_logic ;
  signal GRLFPC2_0_N_124 : std_logic ;
  signal GRLFPC2_0_N_125 : std_logic ;
  signal GRLFPC2_0_N_122 : std_logic ;
  signal GRLFPC2_0_N_96 : std_logic ;
  signal GRLFPC2_0_N_93 : std_logic ;
  signal GRLFPC2_0_N_90 : std_logic ;
  signal GRLFPC2_0_N_64 : std_logic ;
  signal N_12274 : std_logic ;
  signal GRLFPC2_0_RS1V_0_SQMUXA : std_logic ;
  signal N_12275 : std_logic ;
  signal N_12276 : std_logic ;
  signal N_12277 : std_logic ;
  signal N_12278 : std_logic ;
  signal N_12279 : std_logic ;
  signal N_12280 : std_logic ;
  signal N_12281 : std_logic ;
  signal N_12282 : std_logic ;
  signal N_12283 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_592 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_583 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_597 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_580 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_572 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_591 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_593 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_594 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_582 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_600 : std_logic ;
  signal N_12284 : std_logic ;
  signal N_12285 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_613 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_617 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_618 : std_logic ;
  signal N_12286 : std_logic ;
  signal N_12287 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_595 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_587 : std_logic ;
  signal GRLFPC2_0_N_115 : std_logic ;
  signal GRLFPC2_0_N_112 : std_logic ;
  signal GRLFPC2_0_N_111 : std_logic ;
  signal GRLFPC2_0_N_108 : std_logic ;
  signal GRLFPC2_0_N_98 : std_logic ;
  signal GRLFPC2_0_N_83 : std_logic ;
  signal GRLFPC2_0_N_80 : std_logic ;
  signal GRLFPC2_0_N_79 : std_logic ;
  signal GRLFPC2_0_N_76 : std_logic ;
  signal GRLFPC2_0_N_66 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1932 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1933 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_56_I_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_57_I_1 : std_logic ;
  signal GRLFPC2_0_COMB_RS1V_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTRESETORUNIMP : std_logic ;
  signal N_12288 : std_logic ;
  signal N_12289 : std_logic ;
  signal GRLFPC2_0_N_631 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_UN17_INFORCREGSN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN2_NOTDECODEDUNIMP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_7_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_11_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_15_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_17_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_2_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_21_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_25_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_26_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_27_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_32_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_3_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_36_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_37_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_38_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_39_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_40_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_41_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_43_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_45_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_46_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_47_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_50_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_52_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_33_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_34_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_35_I : std_logic ;
  signal GRLFPC2_0_COMB_FPDECODE_ST : std_logic ;
  signal GRLFPC2_0_N_757 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_5_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_54_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_53_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_51_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_49_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_48_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CHECKOVANDDENORM_UN20_NOTPOSSIBLEOV_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CHECKOVANDDENORM_UN20_NOTPOSSIBLEOV_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_UN443_CA_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_57_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN22_GEN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN30_GEN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_UN462_CA_I : std_logic ;
  signal GRLFPC2_0_N_752 : std_logic ;
  signal GRLFPC2_0_N_751 : std_logic ;
  signal N_2362 : std_logic ;
  signal N_8929 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN22_NOTPROP : std_logic ;
  signal GRLFPC2_0_I_237_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_2_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_NE_7 : std_logic ;
  signal GRLFPC2_0_N_636 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_76 : std_logic ;
  signal N_12290 : std_logic ;
  signal N_12291 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_360 : std_logic ;
  signal N_12292 : std_logic ;
  signal N_12293 : std_logic ;
  signal N_12294 : std_logic ;
  signal N_12295 : std_logic ;
  signal N_12296 : std_logic ;
  signal N_12297 : std_logic ;
  signal N_12298 : std_logic ;
  signal N_12299 : std_logic ;
  signal N_12300 : std_logic ;
  signal N_12301 : std_logic ;
  signal N_12302 : std_logic ;
  signal N_12303 : std_logic ;
  signal N_12304 : std_logic ;
  signal N_12305 : std_logic ;
  signal N_12306 : std_logic ;
  signal N_12307 : std_logic ;
  signal N_12308 : std_logic ;
  signal N_12309 : std_logic ;
  signal N_12310 : std_logic ;
  signal N_12311 : std_logic ;
  signal N_12312 : std_logic ;
  signal N_12313 : std_logic ;
  signal N_12314 : std_logic ;
  signal N_12315 : std_logic ;
  signal N_12316 : std_logic ;
  signal N_12317 : std_logic ;
  signal N_12318 : std_logic ;
  signal N_12319 : std_logic ;
  signal N_12320 : std_logic ;
  signal N_12321 : std_logic ;
  signal N_12322 : std_logic ;
  signal N_12323 : std_logic ;
  signal N_12324 : std_logic ;
  signal N_12325 : std_logic ;
  signal N_12326 : std_logic ;
  signal N_12327 : std_logic ;
  signal N_12328 : std_logic ;
  signal N_12329 : std_logic ;
  signal N_12330 : std_logic ;
  signal N_12331 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_11 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_13 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_14 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_15 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_16 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_17 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_19 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_21 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_22 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_23 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_24 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_25 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_27 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_29 : std_logic ;
  signal N_8863 : std_logic ;
  signal N_8825 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_62_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1646 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLOADEN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN4_TOGGLESIG : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN1_TEMP : std_logic ;
  signal GRLFPC2_0_COMB_CCWR4_1 : std_logic ;
  signal GRLFPC2_0_COMB_LOCKGEN_LOCKI_SN_N_10 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_31 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_32 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_36 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_39 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_40 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_41 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_43 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_BUSYMULXFF_UN2_TEMP_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN35_NOTPROP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1880 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1873 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1872 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1871 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1893 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1890 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1888 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1886 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1884 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1883 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1882 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1906 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1904 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1903 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1902 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1897 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1923 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1921 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1899 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1905 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1919 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1920 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1922 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1885 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1891 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1892 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1895 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1874 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1875 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1878 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1924 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1901 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1898 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1896 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1917 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1914 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1915 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1918 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1881 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1909 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1910 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1913 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1912 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1911 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1926 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1916 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1907 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1908 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1900 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1894 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1889 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1887 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1877 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_361 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_STKGEN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN38_GEN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_2 : std_logic ;
  signal GRLFPC2_0_I_237_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW86 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2354 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_EXPBREGLOADEN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLOADEN : std_logic ;
  signal GRLFPC2_0_N_750 : std_logic ;
  signal GRLFPC2_0_COMB_CCWR4 : std_logic ;
  signal GRLFPC2_0_N_737 : std_logic ;
  signal GRLFPC2_0_N_749 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1869 : std_logic ;
  signal GRLFPC2_0_COMB_WRRES4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_45 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_46 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_47 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_49 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_853 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1809 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1808 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_60 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_2 : std_logic ;
  signal N_12332 : std_logic ;
  signal N_12333 : std_logic ;
  signal N_12334 : std_logic ;
  signal N_12335 : std_logic ;
  signal N_12336 : std_logic ;
  signal N_12337 : std_logic ;
  signal N_12338 : std_logic ;
  signal N_12339 : std_logic ;
  signal N_12340 : std_logic ;
  signal N_12341 : std_logic ;
  signal N_12342 : std_logic ;
  signal N_12343 : std_logic ;
  signal N_12344 : std_logic ;
  signal N_12345 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2119 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0 : std_logic ;
  signal GRLFPC2_0_V_FSR_AEXC_1_SQMUXA : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2371 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN20_U_RDN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1748 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1746 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_51 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_54 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_BUSYMULXFF_UN2_TEMP_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN53_GEN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN42_NOTPROP : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_415 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR : std_logic ;
  signal GRLFPC2_0_V_FSR_AEXC_2_SQMUXA : std_logic ;
  signal GRLFPC2_0_V_FSR_CEXC_2_SQMUXA : std_logic ;
  signal GRLFPC2_0_N_797 : std_logic ;
  signal GRLFPC2_0_V_FSR_CEXC_0_SQMUXA : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1741 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_STKGEN_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_35 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_56 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1811 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1810 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1824 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1823 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1820 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1814 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1842 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1840 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1834 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1833 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1831 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1830 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1846 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1845 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1844 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1862 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1816 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1815 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1853 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1839 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1859 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1860 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1861 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1847 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1825 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1826 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1832 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1835 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1865 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1843 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1838 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1837 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1822 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1836 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1812 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1857 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1855 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1858 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1819 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1821 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1850 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1852 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1849 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1851 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1863 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1854 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1856 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1848 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1841 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1829 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1828 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1827 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1818 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1817 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1813 : std_logic ;
  signal N_12346 : std_logic ;
  signal N_12347 : std_logic ;
  signal N_12348 : std_logic ;
  signal N_12349 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_NE_10 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA : std_logic ;
  signal GRLFPC2_0_V_FSR_CEXC_3_SQMUXA : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_800 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1 : std_logic ;
  signal GRLFPC2_0_N_708 : std_logic ;
  signal GRLFPC2_0_COMB_WREN1_9_IV_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_83_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_60_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_95_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_61_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_74_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_59_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_94_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_58_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_109_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_82_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_71_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_87_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_97_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_96_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_84_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_73_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_72_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_81_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_112_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_113_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_110_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_106_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_105_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_101_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_99_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_86_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_85_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_88_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_79_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_108_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_62_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_80_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_65_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_93_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_111_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_67_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_78_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_69_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_98_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_75_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_70_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_90_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_57_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_63_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_89_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_91_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_107_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_92_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_103_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_76_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_104_0 : std_logic ;
  signal N_2376 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_77_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_77_1 : std_logic ;
  signal N_12350 : std_logic ;
  signal N_12351 : std_logic ;
  signal N_12352 : std_logic ;
  signal N_12353 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN49_NOTPROP : std_logic ;
  signal GRLFPC2_0_R_MK_LDOPC_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS : std_logic ;
  signal GRLFPC2_0_N_762 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4 : std_logic ;
  signal N_12354 : std_logic ;
  signal N_12355 : std_logic ;
  signal N_12356 : std_logic ;
  signal N_12357 : std_logic ;
  signal N_12358 : std_logic ;
  signal N_12359 : std_logic ;
  signal N_12360 : std_logic ;
  signal N_12361 : std_logic ;
  signal N_12362 : std_logic ;
  signal N_12363 : std_logic ;
  signal N_12364 : std_logic ;
  signal N_12365 : std_logic ;
  signal N_12366 : std_logic ;
  signal N_12367 : std_logic ;
  signal N_12368 : std_logic ;
  signal N_12369 : std_logic ;
  signal N_12370 : std_logic ;
  signal N_12371 : std_logic ;
  signal N_12372 : std_logic ;
  signal N_12373 : std_logic ;
  signal N_12374 : std_logic ;
  signal N_12375 : std_logic ;
  signal N_12376 : std_logic ;
  signal N_12377 : std_logic ;
  signal N_12378 : std_logic ;
  signal N_12379 : std_logic ;
  signal N_12380 : std_logic ;
  signal N_12381 : std_logic ;
  signal N_12382 : std_logic ;
  signal N_12383 : std_logic ;
  signal N_12384 : std_logic ;
  signal N_12385 : std_logic ;
  signal N_12386 : std_logic ;
  signal N_12387 : std_logic ;
  signal N_12388 : std_logic ;
  signal N_12389 : std_logic ;
  signal N_12390 : std_logic ;
  signal N_12391 : std_logic ;
  signal N_12392 : std_logic ;
  signal N_12393 : std_logic ;
  signal N_12394 : std_logic ;
  signal N_12395 : std_logic ;
  signal N_12396 : std_logic ;
  signal N_12397 : std_logic ;
  signal N_12398 : std_logic ;
  signal N_12399 : std_logic ;
  signal N_12400 : std_logic ;
  signal N_12401 : std_logic ;
  signal N_12402 : std_logic ;
  signal N_12403 : std_logic ;
  signal N_12404 : std_logic ;
  signal N_12405 : std_logic ;
  signal N_12406 : std_logic ;
  signal N_12407 : std_logic ;
  signal N_12408 : std_logic ;
  signal N_12409 : std_logic ;
  signal N_12410 : std_logic ;
  signal N_12411 : std_logic ;
  signal N_12412 : std_logic ;
  signal N_12413 : std_logic ;
  signal N_12414 : std_logic ;
  signal N_12415 : std_logic ;
  signal N_12416 : std_logic ;
  signal N_12417 : std_logic ;
  signal N_12418 : std_logic ;
  signal N_12419 : std_logic ;
  signal N_12420 : std_logic ;
  signal N_12421 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_802 : std_logic ;
  signal N_12422 : std_logic ;
  signal N_12423 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_803 : std_logic ;
  signal N_12424 : std_logic ;
  signal N_12425 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_804 : std_logic ;
  signal N_12426 : std_logic ;
  signal N_12427 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_805 : std_logic ;
  signal N_12428 : std_logic ;
  signal N_12429 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_807 : std_logic ;
  signal N_12430 : std_logic ;
  signal N_12431 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_808 : std_logic ;
  signal N_12432 : std_logic ;
  signal N_12433 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_809 : std_logic ;
  signal N_12434 : std_logic ;
  signal N_12435 : std_logic ;
  signal N_12436 : std_logic ;
  signal N_12437 : std_logic ;
  signal N_12438 : std_logic ;
  signal N_12439 : std_logic ;
  signal N_12440 : std_logic ;
  signal N_12441 : std_logic ;
  signal N_12442 : std_logic ;
  signal N_12443 : std_logic ;
  signal N_12444 : std_logic ;
  signal N_12445 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_806 : std_logic ;
  signal GRLFPC2_0_WREN1_1_SQMUXA_1 : std_logic ;
  signal GRLFPC2_0_N_707 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1743 : std_logic ;
  signal GRLFPC2_0_COMB_FPOP_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1763 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1761 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1760 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1757 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1756 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1755 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1752 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1776 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1774 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1772 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1771 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1766 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1793 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1791 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1789 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1786 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1785 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1781 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1806 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1805 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1802 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1801 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1799 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1796 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1778 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1762 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1769 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1790 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1783 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1782 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1773 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1777 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1779 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1780 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1758 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1795 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1754 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1759 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1768 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1787 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1803 : std_logic ;
  signal N_12446 : std_logic ;
  signal N_12447 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_428 : std_logic ;
  signal N_12448 : std_logic ;
  signal N_12449 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_427 : std_logic ;
  signal N_12450 : std_logic ;
  signal N_12451 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_426 : std_logic ;
  signal N_12452 : std_logic ;
  signal N_12453 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_425 : std_logic ;
  signal N_12454 : std_logic ;
  signal N_12455 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_422 : std_logic ;
  signal N_12456 : std_logic ;
  signal N_12457 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_420 : std_logic ;
  signal N_12458 : std_logic ;
  signal N_12459 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_419 : std_logic ;
  signal N_12460 : std_logic ;
  signal N_12461 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_417 : std_logic ;
  signal N_12462 : std_logic ;
  signal N_12463 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_418 : std_logic ;
  signal N_12464 : std_logic ;
  signal N_12465 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_421 : std_logic ;
  signal N_12466 : std_logic ;
  signal N_12467 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_423 : std_logic ;
  signal N_12468 : std_logic ;
  signal N_12469 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_424 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_344 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN28_STKOUT : std_logic ;
  signal N_12470 : std_logic ;
  signal N_12471 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_459 : std_logic ;
  signal N_12472 : std_logic ;
  signal N_12473 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_462 : std_logic ;
  signal N_12474 : std_logic ;
  signal N_12475 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_465 : std_logic ;
  signal N_12476 : std_logic ;
  signal N_12477 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_479 : std_logic ;
  signal N_12478 : std_logic ;
  signal N_12479 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_483 : std_logic ;
  signal N_12480 : std_logic ;
  signal N_12481 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_487 : std_logic ;
  signal N_12482 : std_logic ;
  signal N_12483 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_493 : std_logic ;
  signal N_12484 : std_logic ;
  signal N_12485 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_495 : std_logic ;
  signal N_12486 : std_logic ;
  signal N_12487 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_489 : std_logic ;
  signal N_12488 : std_logic ;
  signal N_12489 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_448 : std_logic ;
  signal N_12490 : std_logic ;
  signal N_12491 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_492 : std_logic ;
  signal N_12492 : std_logic ;
  signal N_12493 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_460 : std_logic ;
  signal N_12494 : std_logic ;
  signal N_12495 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_470 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1529 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1724 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_506 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_508 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_509 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_510 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_511 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_513 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_514 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_515 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_516 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_517 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_525 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_526 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_528 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_530 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_536 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_539 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_541 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_543 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_544 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_545 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_547 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_549 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_550 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_555 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_556 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_749 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_532 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_523 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_537 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_520 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_512 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_531 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_533 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_534 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_522 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_540 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_553 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_557 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_558 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_535 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_527 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_55_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_0_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_40_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_54_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_35_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_41_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_52_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_39_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_42_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_36_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_19_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_38_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_46_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_44_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_43_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_14_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_13_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_12_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_11_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_10_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_9_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_8_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_49_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_6_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_5_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_3_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_0_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_18_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_32_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_31_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_30_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_29_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_28_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_27_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_26_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_25_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_48_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_20_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_17_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1 : std_logic ;
  signal N_12496 : std_logic ;
  signal N_12497 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_623 : std_logic ;
  signal N_12498 : std_logic ;
  signal N_12499 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_625 : std_logic ;
  signal N_12500 : std_logic ;
  signal N_12501 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_638 : std_logic ;
  signal N_12502 : std_logic ;
  signal N_12503 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_641 : std_logic ;
  signal N_12504 : std_logic ;
  signal N_12505 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_644 : std_logic ;
  signal N_12506 : std_logic ;
  signal N_12507 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_658 : std_logic ;
  signal N_12508 : std_logic ;
  signal N_12509 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_662 : std_logic ;
  signal N_12510 : std_logic ;
  signal N_12511 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_666 : std_logic ;
  signal N_12512 : std_logic ;
  signal N_12513 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_672 : std_logic ;
  signal N_12514 : std_logic ;
  signal N_12515 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_674 : std_logic ;
  signal N_12516 : std_logic ;
  signal N_12517 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_679 : std_logic ;
  signal N_12518 : std_logic ;
  signal N_12519 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_680 : std_logic ;
  signal N_12520 : std_logic ;
  signal N_12521 : std_logic ;
  signal N_12522 : std_logic ;
  signal N_12523 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_624 : std_logic ;
  signal N_12524 : std_logic ;
  signal N_12525 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_668 : std_logic ;
  signal N_12526 : std_logic ;
  signal N_12527 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_627 : std_logic ;
  signal N_12528 : std_logic ;
  signal N_12529 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_671 : std_logic ;
  signal N_12530 : std_logic ;
  signal N_12531 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_639 : std_logic ;
  signal N_12532 : std_logic ;
  signal N_12533 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_649 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_54_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_52_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_39_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_36_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_16_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_15_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_49_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_4_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_1_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_22_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_7_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_29_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_27_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_26_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_25_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_24_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_23_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_48_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_21_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_55_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_2_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_40_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_40_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_54_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_54_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_53_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_51_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_50_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_50_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_50_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_50_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_35_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_35_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_35_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_35_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_41_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_41_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_41_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_52_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_52_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_39_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_39_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_39_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_42_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_42_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_42_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_37_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_37_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_37_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_37_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_36_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_36_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_36_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_19_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_19_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_19_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_38_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_38_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_38_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_46_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_46_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_46_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_45_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_45_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_45_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_45_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_44_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_44_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_44_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_43_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_43_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_43_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_43_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_16_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_16_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_16_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_15_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_15_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_15_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_14_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_14_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_14_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_13_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_13_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_13_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_12_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_12_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_12_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_12_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_11_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_11_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_11_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_10_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_10_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_10_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_10_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_9_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_8_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_47_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_49_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_49_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_49_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_6_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_6_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_34_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_34_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_34_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_34_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_33_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_33_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_33_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_33_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_5_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_5_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_4_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_3_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_2_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_1_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_0_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_0_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_0_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_22_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_22_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_18_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_18_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_18_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_7_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_32_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_32_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_32_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_32_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_31_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_31_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_31_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_31_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_30_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_30_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_29_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_29_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_29_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_28_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_28_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_28_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_27_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_27_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_27_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_26_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_26_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_26_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_25_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_25_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_25_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_24_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_24_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_23_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_23_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_48_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_48_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_21_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_21_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_20_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_20_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_20_4 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_17_2 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_17_3 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_17_4 : std_logic ;
  signal N_12534 : std_logic ;
  signal N_12535 : std_logic ;
  signal N_12536 : std_logic ;
  signal N_12537 : std_logic ;
  signal N_12538 : std_logic ;
  signal N_12539 : std_logic ;
  signal N_12540 : std_logic ;
  signal N_12541 : std_logic ;
  signal N_12542 : std_logic ;
  signal N_12543 : std_logic ;
  signal N_12544 : std_logic ;
  signal N_12545 : std_logic ;
  signal N_12546 : std_logic ;
  signal N_12547 : std_logic ;
  signal N_12548 : std_logic ;
  signal N_12549 : std_logic ;
  signal N_12550 : std_logic ;
  signal N_12551 : std_logic ;
  signal N_12552 : std_logic ;
  signal N_12553 : std_logic ;
  signal N_12554 : std_logic ;
  signal N_12555 : std_logic ;
  signal N_12556 : std_logic ;
  signal N_12557 : std_logic ;
  signal N_12558 : std_logic ;
  signal N_12559 : std_logic ;
  signal N_12560 : std_logic ;
  signal N_12561 : std_logic ;
  signal N_12562 : std_logic ;
  signal N_12563 : std_logic ;
  signal N_12564 : std_logic ;
  signal N_12565 : std_logic ;
  signal N_12566 : std_logic ;
  signal N_12567 : std_logic ;
  signal N_12568 : std_logic ;
  signal N_12569 : std_logic ;
  signal N_12570 : std_logic ;
  signal N_12571 : std_logic ;
  signal N_12572 : std_logic ;
  signal N_12573 : std_logic ;
  signal N_12574 : std_logic ;
  signal N_12575 : std_logic ;
  signal N_12576 : std_logic ;
  signal N_12577 : std_logic ;
  signal N_12578 : std_logic ;
  signal N_12579 : std_logic ;
  signal N_12580 : std_logic ;
  signal N_12581 : std_logic ;
  signal N_12582 : std_logic ;
  signal N_12583 : std_logic ;
  signal N_12584 : std_logic ;
  signal N_12585 : std_logic ;
  signal N_12586 : std_logic ;
  signal N_12587 : std_logic ;
  signal N_12588 : std_logic ;
  signal N_12589 : std_logic ;
  signal N_12590 : std_logic ;
  signal N_12591 : std_logic ;
  signal N_12592 : std_logic ;
  signal N_12593 : std_logic ;
  signal N_12594 : std_logic ;
  signal N_12595 : std_logic ;
  signal N_12596 : std_logic ;
  signal N_12597 : std_logic ;
  signal N_12598 : std_logic ;
  signal N_12599 : std_logic ;
  signal N_12600 : std_logic ;
  signal N_12601 : std_logic ;
  signal N_12602 : std_logic ;
  signal N_12603 : std_logic ;
  signal N_12604 : std_logic ;
  signal N_12605 : std_logic ;
  signal N_12606 : std_logic ;
  signal N_12607 : std_logic ;
  signal N_12608 : std_logic ;
  signal N_12609 : std_logic ;
  signal N_12610 : std_logic ;
  signal N_12611 : std_logic ;
  signal N_12612 : std_logic ;
  signal N_12613 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_40_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_54_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_50_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_50_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_35_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_35_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_41_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_41_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_52_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_39_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_39_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_42_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_42_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_37_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_37_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_36_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_36_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_19_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_19_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_38_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_38_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_46_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_46_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_45_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_45_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_44_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_44_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_43_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_43_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_16_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_16_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_15_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_15_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_14_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_14_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_13_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_13_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_12_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_12_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_11_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_11_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_10_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_10_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_9_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_8_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_49_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_49_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_6_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_34_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_34_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_33_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_33_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_5_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_4_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_3_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_2_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_1_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_0_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_0_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_22_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_18_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_18_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_7_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_32_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_32_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_31_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_31_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_30_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_29_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_29_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_28_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_28_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_27_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_27_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_26_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_26_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_25_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_25_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_24_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_48_5 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_20_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_20_7 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_17_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_17_7 : std_logic ;
  signal N_12614 : std_logic ;
  signal N_12615 : std_logic ;
  signal N_12164 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1519 : std_logic ;
  signal GRLFPC2_0_R_MK_RSTC_1_0 : std_logic ;
  signal GRLFPC2_0_COMB_V_E_AFQ_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_E_AFSR_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_E_FPOP_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_E_LD_1 : std_logic ;
  signal GRLFPC2_0_R_E_AFQ : std_logic ;
  signal GRLFPC2_0_COMB_V_M_AFQ_1 : std_logic ;
  signal GRLFPC2_0_R_E_AFSR : std_logic ;
  signal GRLFPC2_0_COMB_V_M_AFSR_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_M_FPOP_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_M_LD_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1999_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1998_I : std_logic ;
  signal GRLFPC2_0_MOV_5_SQMUXA : std_logic ;
  signal GRLFPC2_0_N_692 : std_logic ;
  signal GRLFPC2_0_COMB_V_FSR_NONSTD_1 : std_logic ;
  signal GRLFPC2_0_N_718_I : std_logic ;
  signal GRLFPC2_0_N_703 : std_logic ;
  signal GRLFPC2_0_N_654 : std_logic ;
  signal GRLFPC2_0_N_657_I : std_logic ;
  signal GRLFPC2_0_N_721_I : std_logic ;
  signal GRLFPC2_0_N_720_I : std_logic ;
  signal GRLFPC2_0_N_637 : std_logic ;
  signal GRLFPC2_0_N_615 : std_logic ;
  signal GRLFPC2_0_N_602 : std_logic ;
  signal GRLFPC2_0_N_728_I : std_logic ;
  signal GRLFPC2_0_N_729_I : std_logic ;
  signal GRLFPC2_0_N_730_I : std_logic ;
  signal GRLFPC2_0_N_731_I : std_logic ;
  signal GRLFPC2_0_N_732_I : std_logic ;
  signal GRLFPC2_0_COMB_V_A_AFQ_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_A_LD_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_A_ST_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_A_AFSR_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_A_SEQERR_1 : std_logic ;
  signal GRLFPC2_0_COMB_RDD_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_372 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1766_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1765_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1764_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1763_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1762_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1761_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1760_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1759_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1758_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1757_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1756_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1755_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1754_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1753_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1752_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1781_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1780_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1779_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1778_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1777_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1776_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1775_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1774_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1773_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1772_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1771_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1770_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1769_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1768_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1767_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1796_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1795_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1794_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1793_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1792_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1791_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1790_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1789_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1788_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1787_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1786_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1785_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1784_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1783_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1782_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1724_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1751_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1806_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1805_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1803_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1802_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1801_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1800_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1799_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1798_I : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1797_I : std_logic ;
  signal GRLFPC2_0_COMB_V_FSR_N_727_I_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_FSR_N_726_I_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_FSR_N_725_I_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_FSR_N_724_I_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_FSR_N_723_I_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_40_I_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_9_6_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_25_0_0_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_33_1_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_34_1_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_47_1_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_47_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_45_1_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_37_1_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_50_1_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_IV_I_141_223_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_35_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_NOTPROP_1_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN30_LOCOV_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN1_S_14_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN20_LOCOV_5_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN20_LOCOV_5 : std_logic ;
  signal G2_2 : std_logic ;
  signal N_12635 : std_logic ;
  signal N_12636 : std_logic ;
  signal G2_4 : std_logic ;
  signal N_12633 : std_logic ;
  signal N_12634 : std_logic ;
  signal G4_2 : std_logic ;
  signal G4_5 : std_logic ;
  signal GRLFPC2_0_R_X_SEQERR_0_0_N_6 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_FAST : std_logic ;
  signal N_12791 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA_1_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_1 : std_logic ;
  signal G0_RN_0 : std_logic ;
  signal G0_SN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1_1 : std_logic ;
  signal N_12941 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_371 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA_M1_E_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_3_1 : std_logic ;
  signal N_12973 : std_logic ;
  signal N_13005 : std_logic ;
  signal N_13009 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_26_0_0X : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_26_0_0_RN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_26_0_0_RN_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_26_0_0_SN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_109 : std_logic ;
  signal N_13011 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA_1 : std_logic ;
  signal N_13062 : std_logic ;
  signal N_13060 : std_logic ;
  signal N_13061 : std_logic ;
  signal N_13088 : std_logic ;
  signal N_13113 : std_logic ;
  signal N_13133 : std_logic ;
  signal N_13154 : std_logic ;
  signal N_13175 : std_logic ;
  signal N_13196 : std_logic ;
  signal N_13217 : std_logic ;
  signal N_13238 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_3 : std_logic ;
  signal N_13323 : std_logic ;
  signal N_13349 : std_logic ;
  signal N_13359 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV_6_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_25_0_0_L9_L7_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_53_I_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_51_I_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_I_SX : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_6_1 : std_logic ;
  signal N_13799 : std_logic ;
  signal N_14071 : std_logic ;
  signal N_14297 : std_logic ;
  signal N_14349 : std_logic ;
  signal N_14348 : std_logic ;
  signal N_14411 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_RN_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_M3_0_SX : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_I_SX : std_logic ;
  signal N_15046 : std_logic ;
  signal N_15069 : std_logic ;
  signal N_15070 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_RN_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_SN : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_21_I_1_0 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_23_I_1_0 : std_logic ;
  signal N_15368 : std_logic ;
  signal N_15367 : std_logic ;
  signal N_15387 : std_logic ;
  signal N_15388 : std_logic ;
  signal N_15389 : std_logic ;
  signal N_13086 : std_logic ;
  signal N_15386 : std_logic ;
  signal N_15385 : std_logic ;
  signal N_15408 : std_logic ;
  signal N_15409 : std_logic ;
  signal N_15410 : std_logic ;
  signal N_13111 : std_logic ;
  signal N_15407 : std_logic ;
  signal N_15406 : std_logic ;
  signal N_15500 : std_logic ;
  signal N_15501 : std_logic ;
  signal N_15502 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_6_I_1 : std_logic ;
  signal N_15543 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_55_I_1 : std_logic ;
  signal N_15777 : std_logic ;
  signal N_15776 : std_logic ;
  signal N_15775 : std_logic ;
  signal N_15809 : std_logic ;
  signal N_15808 : std_logic ;
  signal N_15807 : std_logic ;
  signal N_15822 : std_logic ;
  signal N_15821 : std_logic ;
  signal N_15820 : std_logic ;
  signal N_15854 : std_logic ;
  signal N_15853 : std_logic ;
  signal N_15852 : std_logic ;
  signal N_15885 : std_logic ;
  signal N_15884 : std_logic ;
  signal N_15883 : std_logic ;
  signal N_15898 : std_logic ;
  signal N_15897 : std_logic ;
  signal N_15896 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_9_I_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_5_I_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_30_I_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_7_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_8_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_9_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_10_1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_11_1 : std_logic ;
  signal N_20103 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_REP1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_0_REP1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_6_REP1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_5_REP1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_3_REP1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_2_REP1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_7_REP1 : std_logic ;
  signal GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_4_REP1 : std_logic ;
  signal GRLFPC2_0_R_M_AFQ : std_logic ;
  signal GRLFPC2_0_R_M_AFSR : std_logic ;
  signal GRLFPC2_0_COMB_V_X_AFQ_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_X_AFSR_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_X_FPOP_1 : std_logic ;
  signal GRLFPC2_0_COMB_V_X_LD_1 : std_logic ;
  signal GRLFPC2_0_N_723_I : std_logic ;
  signal GRLFPC2_0_N_724_I : std_logic ;
  signal GRLFPC2_0_N_725_I : std_logic ;
  signal GRLFPC2_0_N_726_I : std_logic ;
  signal GRLFPC2_0_N_727_I : std_logic ;
  component ROM256X1
    generic(
      INIT : bit_vector
    );
    port(
      A0 : in std_logic;
      A1 : in std_logic;
      A2 : in std_logic;
      A3 : in std_logic;
      A4 : in std_logic;
      A5 : in std_logic;
      A6 : in std_logic;
      A7 : in std_logic;
      O : out std_logic  );
  end component;
begin
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_0x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(0),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1997_I,
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_1x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(1),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_5(1),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_2x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(2),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_4(2),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_3x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(3),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_13(3),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_4x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(4),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_14(4),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_5x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(5),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SCTRL_NEW_1,
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_6x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(6),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_16(6),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_7x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1728_I,
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_10x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1741_I,
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_11x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
      D => CPI_D_INST_I(6),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_12x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(12),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_760,
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_13x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(13),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_752,
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_14x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(14),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_1_I(0),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_15x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(15),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_I(42),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_16x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(16),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_RESVEC(0),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_64x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(64),
      D => GRLFPC2_0_N_774_I,
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_65x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(65),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1723_I,
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_66x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(66),
      D => GRLFPC2_0_FPI_START,
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_68x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(68),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN2_NOTDECODEDUNIMP_I,
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_70x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(70),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(68),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_71x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(71),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_UN72_PCTRL_NEW_I,
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_72x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(75),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1519_I,
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_73x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(73),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTRESETORUNIMP_I,
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_74x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(74),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_18(74),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_76x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(76),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_UN61_PCTRL_NEW_I,
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_77x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(77),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14(77),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_78x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(78),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT(7),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_79x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(79),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT(6),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_80x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(80),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT(5),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_81x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(81),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT(4),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_82x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(82),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT(3),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_83x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(83),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT(2),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_84x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(84),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT(1),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_85x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(85),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT(0),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_0: MUXCY_L port map (
      DI => NN_1,
      CI => NN_2,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_0_AND,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_1: MUXCY_L port map (
      DI => NN_1,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_0,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_1_AND,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_2: MUXCY_L port map (
      DI => NN_1,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_1,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_2_AND,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_3: MUXCY_L port map (
      DI => NN_1,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_2,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_3_AND,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_4: MUXCY_L port map (
      DI => NN_1,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_3,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_4_AND,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_5: MUXCY_L port map (
      DI => NN_1,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_4,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_5_AND,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_6: MUXCY_L port map (
      DI => NN_1,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_5,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_6_AND,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_7: MUXCY port map (
      DI => NN_1,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_6,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_7_AND,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT);
  x_grlfpc2_0_r_i_v: FDRE port map (
      Q => GRLFPC2_0_R_I_V,
      D => GRLFPC2_0_COMB_V_I_V_1,
      C => clk,
      R => RST_I,
      CE => GRLFPC2_0_V_I_V_3_SQMUXA_I);
  x_grlfpc2_0_r_mk_busy: FDR port map (
      Q => GRLFPC2_0_R_MK_BUSY,
      D => GRLFPC2_0_COMB_V_MK_BUSY_2,
      C => clk,
      R => RST_I);
  x_grlfpc2_0_r_mk_busy2: FDR port map (
      Q => GRLFPC2_0_R_MK_BUSY2,
      D => GRLFPC2_0_COMB_V_MK_BUSY2_2,
      C => clk,
      R => RST_I);
  x_grlfpc2_0_r_i_exc_0x: FDRE port map (
      Q => GRLFPC2_0_R_I_EXC(0),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1990_I,
      C => clk,
      R => GRLFPC2_0_COMB_UN2_HOLDN,
      CE => GRLFPC2_0_N_762_I);
  x_grlfpc2_0_r_i_exc_1x: FDRE port map (
      Q => GRLFPC2_0_R_I_EXC(1),
      D => GRLFPC2_0_FPO_EXC(1),
      C => clk,
      R => GRLFPC2_0_COMB_UN2_HOLDN,
      CE => GRLFPC2_0_N_762_I);
  x_grlfpc2_0_r_i_exc_2x: FDRE port map (
      Q => GRLFPC2_0_R_I_EXC(2),
      D => GRLFPC2_0_FPO_EXC(2),
      C => clk,
      R => GRLFPC2_0_COMB_UN2_HOLDN,
      CE => GRLFPC2_0_N_762_I);
  x_grlfpc2_0_r_i_exc_3x: FDRE port map (
      Q => GRLFPC2_0_R_I_EXC(3),
      D => GRLFPC2_0_FPO_EXC(3),
      C => clk,
      R => GRLFPC2_0_COMB_UN2_HOLDN,
      CE => GRLFPC2_0_N_762_I);
  x_grlfpc2_0_r_i_exc_4x: FDRE port map (
      Q => GRLFPC2_0_R_I_EXC(4),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1996_I,
      C => clk,
      R => GRLFPC2_0_COMB_UN2_HOLDN,
      CE => GRLFPC2_0_N_762_I);
  x_grlfpc2_0_r_mk_holdn1: FDS port map (
      Q => GRLFPC2_0_R_MK_HOLDN1,
      D => GRLFPC2_0_R_MK_RST2_I,
      C => clk,
      S => RST_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_cry_0: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(257),
      CI => NN_2,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_0,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_cry_1: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(256),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_0,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_1,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_s_1: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_1,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_0,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_cry_2: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(255),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_1,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_2,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_s_2: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_2,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_1,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_cry_3: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(254),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_2,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_3,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_s_3: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_3,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_2,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_cry_4: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(253),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_3,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_4,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_s_4: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_4,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_3,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_cry_5: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(252),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_4,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_5,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_s_5: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_5,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_4,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_cry_6: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(251),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_5,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_6,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_s_6: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_6,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_5,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_cry_7: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(250),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_6,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_7,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_s_7: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_7,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_6,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_cry_8: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(249),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_7,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_8,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_8);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_s_8: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_8,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_7,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_cry_9: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(248),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_8,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_9,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_9);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_s_9: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_9,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_8,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_cry_10: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(247),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_9,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_10,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_10);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_s_10: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_10,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_9,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_cry_11: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(246),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_10,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_11,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_11);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_s_11: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_11,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_10,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_s_12: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_12,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_CRY_11,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_cry_0: MUXCY_L port map (
      DI => NN_1,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_I,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_0,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_s_0: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_0,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_I,
      O => N_2456);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_cry_1: MUXCY_L port map (
      DI => NN_1,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_0,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_1,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_s_1: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_1,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_0,
      O => N_2457);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_cry_2: MUXCY_L port map (
      DI => NN_1,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_1,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_2,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_s_2: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_2,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_1,
      O => N_2458);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_cry_3: MUXCY_L port map (
      DI => NN_1,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_2,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_3,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_s_3: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_3,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_2,
      O => N_2459);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_cry_4: MUXCY_L port map (
      DI => NN_1,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_3,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_4,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_s_4: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_4,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_3,
      O => N_2460);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_cry_5: MUXCY_L port map (
      DI => NN_1,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_4,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_5,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_s_5: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_5,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_4,
      O => N_2461);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_cry_6: MUXCY_L port map (
      DI => NN_1,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_5,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_6,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_s_6: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_6,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_5,
      O => N_2462);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_s_7: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_7,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_CRY_6,
      O => N_2463);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_cry_0: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(0),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_MIXOIN(0),
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_0,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_s_0: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_0,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_MIXOIN(0),
      O => GRLFPC2_0_FPO_EXP(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_cry_1: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(1),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_0,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_1,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_s_1: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_1,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_0,
      O => GRLFPC2_0_FPO_EXP(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_cry_2: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(2),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_1,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_2,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_s_2: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_2,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_1,
      O => GRLFPC2_0_FPO_EXP(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_cry_3: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(3),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_2,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_3,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_s_3: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_3,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_2,
      O => GRLFPC2_0_FPO_EXP(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_cry_4: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(4),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_3,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_4,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_s_4: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_4,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_3,
      O => GRLFPC2_0_FPO_EXP(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_cry_5: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(5),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_4,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_5,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_s_5: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_5,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_4,
      O => GRLFPC2_0_FPO_EXP(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_cry_6: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(6),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_5,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_6,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_s_6: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_6,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_5,
      O => GRLFPC2_0_FPO_EXP(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_cry_7: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(7),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_6,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_7,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_s_7: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_7,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_6,
      O => GRLFPC2_0_FPO_EXP(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_cry_8: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(8),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_7,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_8,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_8);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_s_8: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_8,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_7,
      O => GRLFPC2_0_FPO_EXP(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_cry_9: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(9),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_8,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_9,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_9);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_s_9: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_9,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_8,
      O => GRLFPC2_0_FPO_EXP(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_cry_10: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_998,
      LO => N_2483);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_cry_10_0: MUXCY_L port map (
      DI => N_2483,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_9,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_10,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_10);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_s_10: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_10,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_9,
      O => GRLFPC2_0_FPO_EXP(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_cry_11: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_999,
      LO => N_2490);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_cry_11_0: MUXCY_L port map (
      DI => N_2490,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_10,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_11,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_11);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_s_11: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_11,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_10,
      O => N_2476);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_s_12: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_12,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_CRY_11,
      O => N_2477);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_0: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(0),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN4_TEMP(0),
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_0,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_0: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_0,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN4_TEMP(0),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_1: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(1),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_0,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_1,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_1: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_1,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_0,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_2: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(2),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_1,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_2,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_2: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_2,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_1,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_3: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(3),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_2,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_3,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_3: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_3,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_2,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_4: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(4),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_3,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_4,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_4: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_4,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_3,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_5: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(5),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_4,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_5,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_5: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_5,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_4,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_6: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(6),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_5,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_6,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_6: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_6,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_5,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_7: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(7),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_6,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_7,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_7: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_7,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_6,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_8: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(8),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_7,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_8,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_8);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_8: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_8,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_7,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_9: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(9),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_8,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_9,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_9);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_9: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_9,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_8,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_10: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(10),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_9,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_10,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_10);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_10: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_10,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_9,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_11: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(11),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_10,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_11,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_11);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_11: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_11,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_10,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_12: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(12),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_11,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_12,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_12);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_12: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_12,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_11,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_13: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(13),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_12,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_13,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_13);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_13: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_13,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_12,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_14: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(14),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_13,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_14,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_14);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_14: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_14,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_13,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_15: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(15),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_14,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_15,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_15);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_15: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_15,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_14,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_16: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(16),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_15,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_16,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_16);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_16: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_16,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_15,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_17: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(17),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_16,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_17,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_17);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_17: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_17,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_16,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_18: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(18),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_17,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_18,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_18);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_18: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_18,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_17,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_19: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(19),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_18,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_19,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_19);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_19: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_19,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_18,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_20: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(20),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_19,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_20,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_20);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_20: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_20,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_19,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_21: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(21),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_20,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_21,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_21);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_21: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_21,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_20,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_22: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(22),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_21,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_22,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_22);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_22: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_22,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_21,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_23: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(23),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_22,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_23,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_23);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_23: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_23,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_22,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_24: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(24),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_23,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_24,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_24);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_24: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_24,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_23,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_25: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(25),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_24,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_25,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_25);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_25: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_25,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_24,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_26: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(26),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_25,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_26,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_26);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_26: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_26,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_25,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_27: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(27),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_26,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_27,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_27);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_27: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_27,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_26,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_28: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(28),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_27,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_28,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_28);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_28: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_28,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_27,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_29: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(29),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_28,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_29,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_29);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_29: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_29,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_28,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_30: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(30),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_29,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_30,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_30);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_30: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_30,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_29,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_31: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(31),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_30,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_31,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_31);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_31: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_31,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_30,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_32: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83),
      LO => N_2564);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_32_0: MUXCY_L port map (
      DI => N_2564,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_31,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_32,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_32);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_32: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_32,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_31,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_33: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(82),
      LO => N_2568);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_33_0: MUXCY_L port map (
      DI => N_2568,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_32,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_33,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_33);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_33: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_33,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_32,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_34: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(81),
      LO => N_2572);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_34_0: MUXCY_L port map (
      DI => N_2572,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_33,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_34,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_34);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_34: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_34,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_33,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_35: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(80),
      LO => N_2576);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_35_0: MUXCY_L port map (
      DI => N_2576,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_34,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_35,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_35);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_35: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_35,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_34,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_36: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(79),
      LO => N_2580);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_36_0: MUXCY_L port map (
      DI => N_2580,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_35,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_36,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_36);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_36: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_36,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_35,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_37: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(78),
      LO => N_2584);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_37_0: MUXCY_L port map (
      DI => N_2584,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_36,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_37,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_37);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_37: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_37,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_36,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_38: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(77),
      LO => N_2588);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_38_0: MUXCY_L port map (
      DI => N_2588,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_37,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_38,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_38);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_38: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_38,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_37,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_39: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76),
      LO => N_2592);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_39_0: MUXCY_L port map (
      DI => N_2592,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_38,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_39,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_39);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_39: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_39,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_38,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_40: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75),
      LO => N_2596);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_40_0: MUXCY_L port map (
      DI => N_2596,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_39,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_40,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_40);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_40: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_40,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_39,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_41: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(74),
      LO => N_2600);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_41_0: MUXCY_L port map (
      DI => N_2600,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_40,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_41,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_41);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_41: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_41,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_40,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_42: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(73),
      LO => N_2604);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_42_0: MUXCY_L port map (
      DI => N_2604,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_41,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_42,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_42);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_42: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_42,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_41,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_43: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(72),
      LO => N_2608);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_43_0: MUXCY_L port map (
      DI => N_2608,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_42,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_43,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_43);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_43: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_43,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_42,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_44: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(71),
      LO => N_2612);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_44_0: MUXCY_L port map (
      DI => N_2612,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_43,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_44,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_44);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_44: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_44,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_43,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_45: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(70),
      LO => N_2616);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_45_0: MUXCY_L port map (
      DI => N_2616,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_44,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_45,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_45);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_45: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_45,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_44,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_46: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(69),
      LO => N_2620);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_46_0: MUXCY_L port map (
      DI => N_2620,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_45,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_46,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_46);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_46: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_46,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_45,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_47: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(68),
      LO => N_2624);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_47_0: MUXCY_L port map (
      DI => N_2624,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_46,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_47,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_47);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_47: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_47,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_46,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_48: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(67),
      LO => N_2628);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_48_0: MUXCY_L port map (
      DI => N_2628,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_47,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_48,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_48);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_48: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_48,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_47,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_49: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
      LO => N_2632);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_49_0: MUXCY_L port map (
      DI => N_2632,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_48,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_49,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_49);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_49: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_49,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_48,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_50: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(65),
      LO => N_2636);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_50_0: MUXCY_L port map (
      DI => N_2636,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_49,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_50,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_50);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_50: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_50,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_49,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_51: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
      LO => N_2640);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_51_0: MUXCY_L port map (
      DI => N_2640,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_50,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_51,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_51);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_51: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_51,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_50,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_52: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(63),
      LO => N_2644);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_52_0: MUXCY_L port map (
      DI => N_2644,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_51,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_52,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_52);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_52: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_52,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_51,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_53: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(62),
      LO => N_2648);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_53_0: MUXCY_L port map (
      DI => N_2648,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_52,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_53,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_53);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_53: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_53,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_52,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_54: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(61),
      LO => N_2652);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_54_0: MUXCY_L port map (
      DI => N_2652,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_53,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_54,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_54);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_54: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_54,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_53,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_55: MUXCY_L port map (
      DI => N_20281,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_54,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_55,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_55);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_55: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_55,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_54,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_56: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(59),
      LO => N_2656);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_56_0: MUXCY_L port map (
      DI => N_2656,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_55,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_56,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_56);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_56: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_56,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_55,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_s_57: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_57,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_CRY_56,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_0: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(0),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN4_TEMP(0),
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_0,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_0: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_0,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN4_TEMP(0),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_1: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(1),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_0,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_1,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_1: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_1,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_0,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_2: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(2),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_1,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_2,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_2: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_2,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_1,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_3: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(3),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_2,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_3,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_3: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_3,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_2,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_4: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(4),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_3,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_4,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_4: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_4,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_3,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_5: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(5),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_4,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_5,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_5: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_5,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_4,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_6: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(6),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_5,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_6,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_6: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_6,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_5,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_7: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(7),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_6,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_7,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_7: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_7,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_6,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_8: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(8),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_7,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_8,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_8);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_8: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_8,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_7,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_9: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(9),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_8,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_9,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_9);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_9: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_9,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_8,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_10: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(10),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_9,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_10,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_10);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_10: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_10,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_9,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_11: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(11),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_10,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_11,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_11);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_11: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_11,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_10,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_12: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(12),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_11,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_12,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_12);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_12: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_12,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_11,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_13: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(13),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_12,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_13,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_13);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_13: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_13,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_12,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_14: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(14),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_13,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_14,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_14);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_14: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_14,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_13,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_15: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(15),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_14,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_15,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_15);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_15: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_15,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_14,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_16: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(16),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_15,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_16,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_16);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_16: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_16,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_15,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_17: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(17),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_16,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_17,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_17);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_17: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_17,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_16,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_18: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(18),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_17,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_18,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_18);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_18: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_18,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_17,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_19: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(19),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_18,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_19,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_19);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_19: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_19,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_18,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_20: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(20),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_19,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_20,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_20);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_20: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_20,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_19,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_21: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(21),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_20,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_21,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_21);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_21: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_21,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_20,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_22: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(22),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_21,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_22,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_22);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_22: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_22,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_21,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_23: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(23),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_22,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_23,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_23);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_23: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_23,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_22,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_24: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(24),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_23,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_24,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_24);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_24: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_24,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_23,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_25: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(25),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_24,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_25,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_25);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_25: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_25,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_24,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_26: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(26),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_25,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_26,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_26);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_26: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_26,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_25,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_27: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(27),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_26,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_27,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_27);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_27: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_27,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_26,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_28: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(28),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_27,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_28,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_28);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_28: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_28,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_27,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_29: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(29),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_28,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_29,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_29);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_29: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_29,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_28,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_30: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(30),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_29,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_30,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_30);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_30: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_30,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_29,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_31: MUXCY_L port map (
      DI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(31),
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_30,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_31,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_31);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_31: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_31,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_30,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_32: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83),
      LO => N_2724);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_32_0: MUXCY_L port map (
      DI => N_2724,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_31,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_32,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_32);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_32: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_32,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_31,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_33: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(82),
      LO => N_2731);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_33_0: MUXCY_L port map (
      DI => N_2731,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_32,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_33,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_33);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_33: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_33,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_32,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_34: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(81),
      LO => N_2738);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_34_0: MUXCY_L port map (
      DI => N_2738,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_33,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_34,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_34);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_34: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_34,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_33,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_35: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(80),
      LO => N_2745);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_35_0: MUXCY_L port map (
      DI => N_2745,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_34,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_35,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_35);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_35: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_35,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_34,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_36: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(79),
      LO => N_2752);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_36_0: MUXCY_L port map (
      DI => N_2752,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_35,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_36,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_36);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_36: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_36,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_35,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_37: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(78),
      LO => N_2759);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_37_0: MUXCY_L port map (
      DI => N_2759,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_36,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_37,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_37);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_37: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_37,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_36,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_38: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(77),
      LO => N_2766);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_38_0: MUXCY_L port map (
      DI => N_2766,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_37,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_38,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_38);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_38: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_38,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_37,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_39: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76),
      LO => N_2773);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_39_0: MUXCY_L port map (
      DI => N_2773,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_38,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_39,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_39);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_39: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_39,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_38,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_40: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75),
      LO => N_2780);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_40_0: MUXCY_L port map (
      DI => N_2780,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_39,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_40,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_40);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_40: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_40,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_39,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_41: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(74),
      LO => N_2787);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_41_0: MUXCY_L port map (
      DI => N_2787,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_40,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_41,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_41);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_41: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_41,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_40,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_42: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(73),
      LO => N_2794);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_42_0: MUXCY_L port map (
      DI => N_2794,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_41,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_42,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_42);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_42: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_42,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_41,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_43: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(72),
      LO => N_2801);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_43_0: MUXCY_L port map (
      DI => N_2801,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_42,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_43,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_43);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_43: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_43,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_42,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_44: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(71),
      LO => N_2808);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_44_0: MUXCY_L port map (
      DI => N_2808,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_43,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_44,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_44);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_44: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_44,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_43,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_45: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(70),
      LO => N_2815);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_45_0: MUXCY_L port map (
      DI => N_2815,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_44,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_45,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_45);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_45: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_45,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_44,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_46: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(69),
      LO => N_2822);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_46_0: MUXCY_L port map (
      DI => N_2822,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_45,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_46,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_46);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_46: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_46,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_45,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_47: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(68),
      LO => N_2829);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_47_0: MUXCY_L port map (
      DI => N_2829,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_46,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_47,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_47);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_47: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_47,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_46,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_48: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(67),
      LO => N_2836);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_48_0: MUXCY_L port map (
      DI => N_2836,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_47,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_48,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_48);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_48: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_48,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_47,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_49: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
      LO => N_2843);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_49_0: MUXCY_L port map (
      DI => N_2843,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_48,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_49,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_49);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_49: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_49,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_48,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_50: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(65),
      LO => N_2850);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_50_0: MUXCY_L port map (
      DI => N_2850,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_49,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_50,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_50);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_50: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_50,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_49,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_51: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
      LO => N_2857);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_51_0: MUXCY_L port map (
      DI => N_2857,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_50,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_51,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_51);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_51: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_51,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_50,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_52: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(63),
      LO => N_2864);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_52_0: MUXCY_L port map (
      DI => N_2864,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_51,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_52,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_52);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_52: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_52,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_51,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_53: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(62),
      LO => N_2871);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_53_0: MUXCY_L port map (
      DI => N_2871,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_52,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_53,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_53);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_53: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_53,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_52,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_54: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(61),
      LO => N_2878);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_54_0: MUXCY_L port map (
      DI => N_2878,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_53,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_54,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_54);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_54: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_54,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_53,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_55: MUXCY_L port map (
      DI => N_20279,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_54,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_55,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_55);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_55: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_55,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_54,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_56: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(59),
      LO => N_2885);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_56_0: MUXCY_L port map (
      DI => N_2885,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_55,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_56,
      LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_56);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_56: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_56,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_55,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_s_57: XORCY port map (
      LI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_57,
      CI => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_CRY_56,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_pctrl_67x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(67),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2032_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_9x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(9),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN20_U_RDN_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1749_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_8x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(8),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1748_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1749_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_374x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(374),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_115_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELECTDIVMULT_UN86_DIVMULTV);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_375x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(375),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_I(375),
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_I(375));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_376x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(376),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2297,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2298);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_245x: FDR port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(245),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_2,
      C => clk,
      R => RST_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_246x: FDR port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(246),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_1,
      C => clk,
      R => RST_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_232x: FDR port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(232),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_814,
      C => clk,
      R => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_815);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_233x: FDR port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(233),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_813,
      C => clk,
      R => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_815);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_234x: FDR port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(234),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_812,
      C => clk,
      R => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_815);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_235x: FDR port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(235),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_811,
      C => clk,
      R => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_815);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_236x: FDR port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(236),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_810,
      C => clk,
      R => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_815);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_162x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(162),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_113_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(162));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_163x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(163),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_112_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(163));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_164x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(164),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_111_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(164));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_165x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(165),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_110_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(165));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_166x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(166),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_109_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(166));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_167x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(167),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_108_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(167));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_168x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(168),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_107_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(168));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_169x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(169),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_106_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(169));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_170x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(170),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_105_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(170));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_171x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(171),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_104_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14_M(171));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_172x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(172),
      D => N_8694_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2342);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_173x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(173),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_102_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(173));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_147x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(147),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_101_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(147));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_148x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(148),
      D => N_8699_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2207);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_149x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(149),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_99_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(149));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_150x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(150),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_98_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(150));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_151x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(151),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_97_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(151));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_152x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(152),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_96_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(152));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_153x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(153),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_95_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(153));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_154x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(154),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_94_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(154));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_155x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(155),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_93_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(155));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_156x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(156),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_92_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(156));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_157x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(157),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_91_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(157));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_158x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(158),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_90_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(158));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_159x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(159),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_89_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(159));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_160x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(160),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_88_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(160));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_161x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(161),
      D => N_8692_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2338);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_132x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(132),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_86_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(132));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_133x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(133),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_85_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(133));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_134x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(134),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_84_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(134));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_135x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(135),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_83_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(135));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_136x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(136),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_82_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(136));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_137x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(137),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_81_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(137));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_138x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(138),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_80_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(138));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_139x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(139),
      D => N_8693_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2323);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_140x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(140),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_78_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(140));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_141x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(141),
      D => N_8688_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2328);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_142x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(142),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_76_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14_M(142));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_143x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(143),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_75_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(143));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_144x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(144),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_74_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(144));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_145x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(145),
      D => N_8689_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2334);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_146x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(146),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_72_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(146));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_117x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(117),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_71_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(117));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_118x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(118),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_70_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(118));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_119x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(119),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_69_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(119));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_120x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(120),
      D => N_8700_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2302);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_121x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(121),
      D => N_8690_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2305);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_122x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(122),
      D => N_8701_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2309);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_123x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(123),
      D => N_8691_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2312);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_124x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(124),
      D => N_8702_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2316);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_125x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(125),
      D => N_8687_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2319);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_126x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(126),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_62_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(126));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_127x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(127),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_61_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(127));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_128x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(128),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_60_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(128));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_129x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(129),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_59_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(129));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_130x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(130),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_58_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(130));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_131x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(131),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_57_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(131));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_115x: FDR port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(115),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_0,
      C => clk,
      R => RST_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_116x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(116),
      D => N_8703_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2299);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_57x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(57),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_55_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_42x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(42),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_54_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_43x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(43),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_53_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_44x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(44),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_52_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_45x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(45),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_51_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_46x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(46),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_50_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_47x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(47),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_49_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_48x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(48),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_48_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_49x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(49),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_47_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_50x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(50),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_46_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_51x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_45_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_52x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(52),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_44_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_53x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_43_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_54x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(54),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_42_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_55x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_41_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_56x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(56),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_40_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0_M(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_27x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(27),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_39_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_28x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(28),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_38_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_29x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(29),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_37_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_30x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(30),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_36_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_31x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(31),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_35_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_32x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(32),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_34_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_33x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(33),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_33_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_34x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(34),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_32_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_35x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(35),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_31_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_36x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(36),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_30_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_37x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(37),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_29_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_38x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(38),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_28_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_39x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(39),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_27_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_40x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(40),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_26_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_41x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(41),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_25_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_12x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(12),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_24_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_13x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(13),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_23_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_14x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(14),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_22_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_15x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(15),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_21_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_16x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(16),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_20_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_17x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_19_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_18x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(18),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_18_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_19x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_17_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_20x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(20),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_16_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_21x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_15_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_22x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(22),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_14_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_23x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_13_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_24x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(24),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_12_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_25x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(25),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_11_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_26x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(26),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_10_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_0x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(0),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_9_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_1x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_8_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_2x: FDR port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(2),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC,
      C => clk,
      R => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0_I_M(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_3x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_7_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_4x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_6_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_5x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_5_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_6x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(6),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_4_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_7x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(7),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_3_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_8x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_2_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_9x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(9),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_1_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_10x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(10),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_0_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_11x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(11),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_I,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(46));
  x_grlfpc2_0_r_mk_ldop: FDR port map (
      Q => GRLFPC2_0_R_MK_LDOP,
      D => GRLFPC2_0_R_MK_LDOPC,
      C => clk,
      R => CPI_D_INST_I(31));
  x_grlfpc2_0_r_mk_rst: FDR port map (
      Q => GRLFPC2_0_R_MK_RST,
      D => GRLFPC2_0_R_MK_RSTC,
      C => clk,
      R => HOLDN_I);
  x_grlfpc2_0_r_a_rs2_0x: FDRE port map (
      Q => GRLFPC2_0_R_A_RS2(0),
      D => cpi_d_inst(0),
      C => clk,
      R => GRLFPC2_0_COMB_RS2_1_SN_N_2,
      CE => holdn);
  x_grlfpc2_0_r_a_rs2_1x: FDRE port map (
      Q => GRLFPC2_0_R_A_RS2(1),
      D => cpi_d_inst(1),
      C => clk,
      R => GRLFPC2_0_COMB_RS2_1_SN_N_2,
      CE => holdn);
  x_grlfpc2_0_r_a_rs2_2x: FDRE port map (
      Q => GRLFPC2_0_R_A_RS2(2),
      D => cpi_d_inst(2),
      C => clk,
      R => GRLFPC2_0_COMB_RS2_1_SN_N_2,
      CE => holdn);
  x_grlfpc2_0_r_a_rs2_3x: FDRE port map (
      Q => GRLFPC2_0_R_A_RS2(3),
      D => cpi_d_inst(3),
      C => clk,
      R => GRLFPC2_0_COMB_RS2_1_SN_N_2,
      CE => holdn);
  x_grlfpc2_0_r_a_rs2_4x: FDRE port map (
      Q => GRLFPC2_0_R_A_RS2(4),
      D => cpi_d_inst(4),
      C => clk,
      R => GRLFPC2_0_COMB_RS2_1_SN_N_2,
      CE => holdn);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_0: ROM256X1 
  generic map(
    INIT => X"083000E400480800020020000000004D08020480300000310000008000002000"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6829_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_1: ROM256X1 
  generic map(
    INIT => X"0000004802A000008A001028000082042848008C0B0000000288088A22AA0000"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6830_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_2: ROM256X1 
  generic map(
    INIT => X"023A02C822E89B3BCECEF77E9999B2DDAC6E66ACEB8B80B1EFDE7DFEBFFBED34"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6831_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_3: ROM256X1 
  generic map(
    INIT => X"0035008822A0111BC216F21C100532542C49228C0B0B008083CA015E26BB4C00"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6832_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_4: ROM256X1 
  generic map(
    INIT => X"0027025832ACB3608645111801588204283E24BC8B8480C84F8E742A37BB8C20"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6833_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_5: ROM256X1 
  generic map(
    INIT => X"002502D832A429488E491116817D921D287840BCAB028079E798444E37EA6014"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6834_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_6: ROM256X1 
  generic map(
    INIT => X"003F001912ACBB6E8E9CB76C004632CDAC4F041DE38F00FDAF86199A26AAA520"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6835_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_7: ROM256X1 
  generic map(
    INIT => X"021D00982004904002CF954009B800D08C60223088098048E10E45389DC84D14"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6836_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_8: ROM256X1 
  generic map(
    INIT => X"021D00D822A41048C68AE2229881A254A41A22BC030D80C8A6D6299AAAAA4510"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6837_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_9: ROM256X1 
  generic map(
    INIT => X"022702C002EC823B8C8595460004A200285E64A4C3848000AED6302222730400"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6838_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_10: ROM256X1 
  generic map(
    INIT => X"022A02C83040221B009EA66688C88094804B62AC8102808081C008C4AE33CD32"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6839_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_11: ROM256X1 
  generic map(
    INIT => X"003402800000082A40026018100020C900032428A80B00B1890000B004006800"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6840_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_12: ROM256X1 
  generic map(
    INIT => X"000000910000084C020000280002000D880220B9210000FD0100080006026800"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6841_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_13: ROM256X1 
  generic map(
    INIT => X"020002110000A86E0088202000020009002204192002007D8910089006402002"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6842_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_14: ROM256X1 
  generic map(
    INIT => X"0230005902E8A844C08A6312100282CDA8640495AA09007D0A08019A2000A822"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6843_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_15: ROM256X1 
  generic map(
    INIT => X"023B00C832ECBB13CED7D75E99FDB2DDAC7C668CEB8D80B1EECE75EEBBBBAD36"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6844_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_16: ROM256X1 
  generic map(
    INIT => X"00000011000000440000000000020000000000110000004C0000000000000000"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6845_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_17: ROM256X1 
  generic map(
    INIT => X"0001001100040044000000000000000000010011000400440000000000000000"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6846_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_18: ROM256X1 
  generic map(
    INIT => X"0000082080000000000000002000002140000000002000008020020000008000"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6847_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_19: ROM256X1 
  generic map(
    INIT => X"0000002000000002000000002000000000000000100200008080000000000000"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6848_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_20: ROM256X1 
  generic map(
    INIT => X"FFFFFFDFFFFFFFFDEFEFFFFFDFFFDFFFEEEEFFFFEBF9FFFD7F7FFFFFFFFFFFFF"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6849_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_21: ROM256X1 
  generic map(
    INIT => X"000013000000440000000080020000000000110000004C000000000000000000"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6850_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_22: ROM256X1 
  generic map(
    INIT => X"FF7FFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFF"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6851_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_23: ROM256X1 
  generic map(
    INIT => X"3080A000400200800000000000000D0202800002000031000000800000000000"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6852_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_24: ROM256X1 
  generic map(
    INIT => X"3080E400080300800000000000000D0202000002000031000000800000000000"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6853_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_25: ROM256X1 
  generic map(
    INIT => X"3080A000480300802000000000000D0202808000000031000000000000000000"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6854_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_26: ROM256X1 
  generic map(
    INIT => X"2A853BB18805EC4C00880089220240294122B9F134204CFFA1A342210400E822"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6855_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_27: ROM256X1 
  generic map(
    INIT => X"0000000000020080000000000000090680000000000031000000000000000150"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6856_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_28: ROM256X1 
  generic map(
    INIT => X"070F131114044F4C20890088020624002221511102144C4C2812400000404802"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6857_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_29: ROM256X1 
  generic map(
    INIT => X"22853BB18115E44401880089264220296123B1B124244CFFA13342210440E822"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6858_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_30: ROM256X1 
  generic map(
    INIT => X"4800082888C02002000109082004422161C228E0143200928BB002222440C022"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6859_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_31: ROM256X1 
  generic map(
    INIT => X"4D0F13191DD66FCE2101098806466F06A3C379F116167DDE0B90002224404172"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6860_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_32: ROM256X1 
  generic map(
    INIT => X"4502000004000A08000000000000000003020020061000820910002004400000"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6861_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_33: ROM256X1 
  generic map(
    INIT => X"0502000804000A0A000000000000000003022020061200820910002004400000"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6862_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_34: ROM256X1 
  generic map(
    INIT => X"00000131000004440004100022920000002001114000044C8000004090010000"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6863_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_35: ROM256X1 
  generic map(
    INIT => X"0F2F091995F42F5F8905110006D62225E16B69B1563604FE2AA2424290030920"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6864_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_36: ROM256X1 
  generic map(
    INIT => X"000000110000804C000400000002000000220031400000CCA302006804810000"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6865_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_37: ROM256X1 
  generic map(
    INIT => X"4000001300C0814C000409000002000000224031400000DDA212004820C10052"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6866_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_38: ROM256X1 
  generic map(
    INIT => X"FFFEFFFFFFFBFFFFBB3FBBBBFFFFFDFFFFFEFFBF6FBBFFFFBB3ABBFFFDFFFFFF"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6867_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_39: ROM256X1 
  generic map(
    INIT => X"0001000000040000444044450000020000010000800400004444440000200000"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6868_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_40: ROM256X1 
  generic map(
    INIT => X"FFFEFFFFFFFBFFFFBB3FBBBBFFFFFDFFFFFEFFFF6FBBFFFFBB3BBBFFFDDFFFFF"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6869_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_41: ROM256X1 
  generic map(
    INIT => X"0000002000000000000000000020000000000000000000008000000000000000"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6870_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_42: ROM256X1 
  generic map(
    INIT => X"0000000000000008000000000000000000020000000200800000000000000000"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6871_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_43: ROM256X1 
  generic map(
    INIT => X"ED4FFFA6E507DD9332B1B8A923443D3EDF9BF3CA75F6FF23B8B3BAB142E87FD7"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6872_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_44: ROM256X1 
  generic map(
    INIT => X"121000000A2000084C4EC6449899C0410024042400010080454C454C9D130000"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6873_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_45: ROM256X1 
  generic map(
    INIT => X"4560005914D820648100011244020280204000118808007D02000002200482AA"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6874_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_46: ROM256X1 
  generic map(
    INIT => X"00002000400200802000000000000D0688808080000031000000000000000000"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6875_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_47: ROM256X1 
  generic map(
    INIT => X"FF7FFFFFCFFFDFDFFFFFFFFFFFFFFFF7FFF7F7FFFFFFFFFFFFFFFFFFFFFBDF77"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6876_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_48: ROM256X1 
  generic map(
    INIT => X"0005000000041100000000000000100000004000000000000000000000000080"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6877_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_49: ROM256X1 
  generic map(
    INIT => X"2010805112212A644002C20110228048020400552201007D1009010940042008"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6878_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_50: ROM256X1 
  generic map(
    INIT => X"0520000804C80000810001120400028020400000880800000200000220000800"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6879_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_51: ROM256X1 
  generic map(
    INIT => X"3FB580593FFD3B6CCD4EC757DCFBD2C9226C4C75AA1900FD5F5D454FFD57A8A8"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6880_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_52: ROM256X1 
  generic map(
    INIT => X"00002000400200802000000000000D0688808080000031000000000000000000"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6881_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_53: ROM256X1 
  generic map(
    INIT => X"4040000000000000000000000000000000000000000000000000000000000202"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6882_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_54: ROM256X1 
  generic map(
    INIT => X"404000001000202000000000000000000000000000000000000000000004020A"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6883_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_55: ROM256X1 
  generic map(
    INIT => X"00001B208000440210100080220020215111110014264E1290A0020040008020"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6884_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_56: ROM256X1 
  generic map(
    INIT => X"05051BB1970475665055548032D6302151115311142E4E4EE0A6531490058008"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6885_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_57: ROM256X1 
  generic map(
    INIT => X"0800000831C82A20080081100060020820480800801002311A00000240062008"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6886_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_58: ROM256X1 
  generic map(
    INIT => X"4545001915DCA06E400545105046020000600031800A00CC220601140005020A"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6887_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_59: ROM256X1 
  generic map(
    INIT => X"4040000011103120000000004040100000004000000000000010000020440A8A"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6888_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_60: ROM256X1 
  generic map(
    INIT => X"4045000000040000010000000400000000000000000000000000000000000202"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6889_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_61: ROM256X1 
  generic map(
    INIT => X"454000001510202000000000404000000000000000000000000000000004020A"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6890_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_00_62: ROM256X1 
  generic map(
    INIT => X"0705000004040008044C0444889920000021042000040080454444449D110008"
  )
  port map (
    A0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
    A1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
    A2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
    A3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
    A4 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
    A5 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
    A6 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
    A7 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
    O => N_6891_A);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_53x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(62),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expybus_2_6x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(30),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPYBUS_2(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m5s2: LUT2 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(11),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(12),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SM3_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_stickyforsr1: LUT2 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(56),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(57),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2030);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_RomxzSL2FromC: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_ROMXZSL2FROMC);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_7_and1: LUT2 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(54),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_7_AND1);
  x_grlfpc2_0_fpco_holdn: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_R_MK_HOLDN1,
    I1 => GRLFPC2_0_R_MK_HOLDN2,
    O => cpo_holdn);
  x_grlfpc2_0_comb_un10_iuexec: LUT2 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => GRLFPC2_0_R_MK_RST,
    I1 => GRLFPC2_0_R_MK_RST2,
    O => GRLFPC2_0_N_782);
  x_grlfpc2_0_comb_pexc9: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_R_STATE(0),
    I1 => GRLFPC2_0_R_STATE(1),
    O => CPO_EXC_INT_2);
  x_grlfpc2_0_comb_qne2: LUT2 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => GRLFPC2_0_R_STATE(0),
    I1 => GRLFPC2_0_R_STATE(1),
    O => GRLFPC2_0_SEQERR_1_SQMUXA_1_SN);
  x_grlfpc2_0_mov_0_sqmuxa_2: LUT2 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => cpi_d_inst(10),
    I1 => cpi_d_inst(11),
    O => GRLFPC2_0_MOV_0_SQMUXA_2);
  x_grlfpc2_0_mov_2_sqmuxa_2: LUT2 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => cpi_d_inst(11),
    I1 => cpi_d_inst(12),
    O => GRLFPC2_0_MOV_2_SQMUXA_2);
  x_grlfpc2_0_comb_fpdecode_mov6_2: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => cpi_d_inst(11),
    I1 => cpi_d_inst(12),
    O => GRLFPC2_0_COMB_FPDECODE_MOV6_2);
  x_grlfpc2_0_comb_fpdecode_afq12: LUT2 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => cpi_d_inst(30),
    I1 => cpi_d_inst(31),
    O => GRLFPC2_0_COMB_FPDECODE_AFQ12);
  x_grlfpc2_0_comb_fpdecode_afq13: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => cpi_d_inst(30),
    I1 => cpi_d_inst(31),
    O => GRLFPC2_0_COMB_FPDECODE_AFQ13);
  x_grlfpc2_0_comb_v_e_stdata2: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => cpi_a_cnt(0),
    I1 => cpi_a_cnt(1),
    O => GRLFPC2_0_COMB_V_E_STDATA2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_2x: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(371),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_0x: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(373),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_17x: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(356),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(17));
  x_grlfpc2_0_comb_un22_ccv: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => cpi_m_inst(19),
    I1 => GRLFPC2_0_R_M_FPOP,
    O => GRLFPC2_0_COMB_UN22_CCV);
  x_grlfpc2_0_comb_un14_ccv: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => cpi_x_inst(19),
    I1 => GRLFPC2_0_R_X_FPOP,
    O => GRLFPC2_0_COMB_UN14_CCV);
  x_grlfpc2_0_annulres_0_sqmuxa_3_2: LUT2 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => GRLFPC2_0_R_E_FPOP,
    I1 => GRLFPC2_0_R_M_FPOP,
    O => GRLFPC2_0_ANNULRES_0_SQMUXA_3_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_36x: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(337),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_40x: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(333),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_sftlft_aregxorbreg: LUT2 
  generic map(
    INIT => X"6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(12),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(13),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_AREGXORBREG);
  x_grlfpc2_0_v_fsr_nonstd_0_sqmuxa: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_R_X_AFSR,
    I1 => GRLFPC2_0_R_X_LD,
    O => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA);
  x_grlfpc2_0_comb_wren22: LUT2 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => cpi_x_cnt(0),
    I1 => cpi_x_cnt(1),
    O => GRLFPC2_0_COMB_WREN22);
  x_grlfpc2_0_comb_mexc_1_4x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_R_FSR_TEM(4),
    I1 => GRLFPC2_0_R_I_EXC(4),
    O => GRLFPC2_0_COMB_MEXC_1(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_sftlft_un1_grfpus: LUT2 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(65),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_I(24),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2031);
  x_grlfpc2_0_I_237_1: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => cpi_d_inst(21),
    I1 => cpi_d_inst(24),
    O => GRLFPC2_0_N_703_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m8s2: LUT2 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(7),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SM6_I);
  x_grlfpc2_0_mov_2_sqmuxa_1_0: LUT2 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => cpi_d_inst(5),
    I1 => cpi_d_inst(6),
    O => GRLFPC2_0_MOV_2_SQMUXA_1_0);
  x_grlfpc2_0_mov_0_sqmuxa_3: LUT2 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => cpi_d_inst(7),
    I1 => cpi_d_inst(8),
    O => GRLFPC2_0_MOV_0_SQMUXA_3);
  x_grlfpc2_0_comb_mexc_1_3x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_R_FSR_TEM(3),
    I1 => GRLFPC2_0_R_I_EXC(3),
    O => GRLFPC2_0_COMB_MEXC_1(3));
  x_grlfpc2_0_comb_mexc_1_2x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_R_FSR_TEM(2),
    I1 => GRLFPC2_0_R_I_EXC(2),
    O => GRLFPC2_0_COMB_MEXC_1(2));
  x_grlfpc2_0_comb_mexc_1_1x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_R_FSR_TEM(1),
    I1 => GRLFPC2_0_R_I_EXC(1),
    O => GRLFPC2_0_COMB_MEXC_1(1));
  x_grlfpc2_0_comb_mexc_1_0x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_R_FSR_TEM(0),
    I1 => GRLFPC2_0_R_I_EXC(0),
    O => GRLFPC2_0_COMB_MEXC_1(0));
  x_grlfpc2_0_comb_un1_fpci_1: LUT2 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => cpi_m_annul,
    I1 => cpi_m_trap,
    O => GRLFPC2_0_COMB_UN1_FPCI_1_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_t_3_i_o2_0_0x: LUT2 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(374),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(376),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2281_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_entryshft_s_3: LUT2 
  generic map(
    INIT => X"6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(80),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(81),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_ENTRYSHFT_S_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_feedbackmulxff_un19_feedback_2: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(51),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(52),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN19_FEEDBACK_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m2s2: LUT2 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(15),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(16),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SM0_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_lib_0x: LUT2 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(10),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(44),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_LIB(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_55x: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(318),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_42x: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(331),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_37x: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(336),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_26x: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(347),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_2_30x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_16_REP1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un23_temp: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(74),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(75),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN23_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un2_temp: LUT2 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(75),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(76),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_temp: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(42),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(15),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_conditional_6x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(9),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_CONDITIONAL(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_axb_0: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(244),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(257),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_axb_12: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(232),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(245),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_12);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_axb_7: LUT1 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(78),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_r_dpath_inv_4_0: LUT2 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(13),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(14),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV_4_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un5_notshiftcount1_0: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(14),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(16),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN5_NOTSHIFTCOUNT1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_r_sctrl_2_sn_m1_e_0: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(25),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(26),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_2_SN_M1_E_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_mixoin_0_0x: LUT3 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(35),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_MIXOIN(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un1_waitq_0_0x: LUT3 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(58),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_I(19),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_55x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(60),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(18),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_topbitsin_0_0x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(244),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(44),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_topbitsin_0_1x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(243),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(44),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_topbitsin_0_3x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(241),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(44),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_topbitsin_0_4x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(240),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(44),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_topbitsin_0_5x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(239),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(44),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_topbitsin_0_7x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(237),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(44),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_topbitsin_0_8x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(44),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(12),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_0_0x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(25),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(57),
    I2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_0_1x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(24),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(56),
    I2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_0_2x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_0_3x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(22),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(54),
    I2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_0_4x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_0_5x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(20),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(52),
    I2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_0_6x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_0_7x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(18),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(50),
    I2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notmultip_0_8x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(49),
    I2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_2_0_4x: LUT3_L 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(240),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(253),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_992);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_2_0_10x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(234),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(247),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_998);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_2_0_11x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(233),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(246),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_999);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_2_0_12x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(232),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(245),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1000);
  x_grlfpc2_0_comb_dbgdata_5_0_0_0x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => rfo1_data1(0),
    I2 => rfo2_data1(0),
    O => GRLFPC2_0_N_311);
  x_grlfpc2_0_comb_dbgdata_5_0_0_1x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => rfo1_data1(1),
    I2 => rfo2_data1(1),
    O => GRLFPC2_0_N_312);
  x_grlfpc2_0_comb_dbgdata_5_0_0_2x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => rfo1_data1(2),
    I2 => rfo2_data1(2),
    O => GRLFPC2_0_N_313);
  x_grlfpc2_0_comb_dbgdata_5_0_0_3x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => rfo1_data1(3),
    I2 => rfo2_data1(3),
    O => GRLFPC2_0_N_314);
  x_grlfpc2_0_comb_dbgdata_5_0_0_5x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => rfo1_data1(5),
    I2 => rfo2_data1(5),
    O => GRLFPC2_0_N_316);
  x_grlfpc2_0_comb_dbgdata_5_0_0_6x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => rfo1_data1(6),
    I2 => rfo2_data1(6),
    O => GRLFPC2_0_N_317);
  x_grlfpc2_0_comb_dbgdata_5_0_0_7x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => rfo1_data1(7),
    I2 => rfo2_data1(7),
    O => GRLFPC2_0_N_318);
  x_grlfpc2_0_comb_dbgdata_5_0_0_8x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => rfo1_data1(8),
    I2 => rfo2_data1(8),
    O => GRLFPC2_0_N_319);
  x_grlfpc2_0_comb_dbgdata_5_0_0_9x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => rfo1_data1(9),
    I2 => rfo2_data1(9),
    O => GRLFPC2_0_N_320);
  x_grlfpc2_0_comb_dbgdata_5_0_0_10x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => rfo1_data1(10),
    I2 => rfo2_data1(10),
    O => GRLFPC2_0_N_321);
  x_grlfpc2_0_comb_dbgdata_5_0_0_11x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => rfo1_data1(11),
    I2 => rfo2_data1(11),
    O => GRLFPC2_0_N_322);
  x_grlfpc2_0_comb_dbgdata_5_0_0_22x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => rfo1_data1(22),
    I2 => rfo2_data1(22),
    O => GRLFPC2_0_N_333);
  x_grlfpc2_0_comb_dbgdata_5_0_0_23x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => rfo1_data1(23),
    I2 => rfo2_data1(23),
    O => GRLFPC2_0_N_334);
  x_grlfpc2_0_comb_dbgdata_5_0_0_24x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => rfo1_data1(24),
    I2 => rfo2_data1(24),
    O => GRLFPC2_0_N_335);
  x_grlfpc2_0_comb_dbgdata_5_0_0_25x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => rfo1_data1(25),
    I2 => rfo2_data1(25),
    O => GRLFPC2_0_N_336);
  x_grlfpc2_0_comb_dbgdata_5_0_0_27x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => rfo1_data1(27),
    I2 => rfo2_data1(27),
    O => GRLFPC2_0_N_338);
  x_grlfpc2_0_comb_dbgdata_5_0_0_30x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => rfo1_data1(30),
    I2 => rfo2_data1(30),
    O => GRLFPC2_0_N_341);
  x_grlfpc2_0_comb_dbgdata_5_0_0_31x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => rfo1_data1(31),
    I2 => rfo2_data1(31),
    O => GRLFPC2_0_N_342);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_topbitsin_0_2x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(242),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(44),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(2));
  x_grlfpc2_0_comb_dbgdata_5_0_0_14x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => rfo1_data1(14),
    I2 => rfo2_data1(14),
    O => GRLFPC2_0_N_325);
  x_grlfpc2_0_comb_dbgdata_5_0_0_4x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => rfo1_data1(4),
    I2 => rfo2_data1(4),
    O => GRLFPC2_0_N_315);
  x_grlfpc2_0_comb_dbgdata_5_0_0_26x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => rfo1_data1(26),
    I2 => rfo2_data1(26),
    O => GRLFPC2_0_N_337);
  x_grlfpc2_0_comb_dbgdata_5_0_0_16x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => rfo1_data1(16),
    I2 => rfo2_data1(16),
    O => GRLFPC2_0_N_327);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_topbitsin_0_6x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(238),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(44),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_SelInitRemBit: LUT3 
  generic map(
    INIT => X"04"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(5),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELINITREMBIT);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_expybus_1_3x: LUT3 
  generic map(
    INIT => X"51"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2017);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_expybus_1_1x: LUT3_L 
  generic map(
    INIT => X"15"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP1,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2016);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_computeconst_un49_resvec: LUT3 
  generic map(
    INIT => X"40"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_COMPUTECONST_UN49_RESVEC);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_notam2_0: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2030,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_NOTAM2_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_feedbackmulxff_un19_feedback: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN19_FEEDBACK_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(49),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(50),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN19_FEEDBACK);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_sftlft_un5_temp: LUT3 
  generic map(
    INIT => X"07"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(27),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(28),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(65),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_3_SN_I3_I_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_status_1_6x: LUT3 
  generic map(
    INIT => X"5D"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(38),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(40),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2003);
  x_grlfpc2_0_comb_un1_r_i_v: LUT3 
  generic map(
    INIT => X"40"
  )
  port map (
    I0 => GRLFPC2_0_R_I_EXEC,
    I1 => GRLFPC2_0_R_I_V,
    I2 => GRLFPC2_0_R_X_FPOP,
    O => GRLFPC2_0_COMB_UN1_R_I_V);
  x_grlfpc2_0_comb_fpdecode_afq5_2: LUT3 
  generic map(
    INIT => X"10"
  )
  port map (
    I0 => cpi_d_inst(22),
    I1 => cpi_d_inst(23),
    I2 => GRLFPC2_0_N_703_1,
    O => GRLFPC2_0_COMB_FPDECODE_AFQ4_1);
  x_grlfpc2_0_comb_fpdecode_afq7_1: LUT4 
  generic map(
    INIT => X"0100"
  )
  port map (
    I0 => cpi_d_inst(21),
    I1 => cpi_d_inst(22),
    I2 => cpi_d_inst(23),
    I3 => cpi_d_inst(24),
    O => GRLFPC2_0_COMB_FPDECODE_AFQ7_1);
  x_grlfpc2_0_comb_fpdecode_afq2_2: LUT3 
  generic map(
    INIT => X"10"
  )
  port map (
    I0 => cpi_d_inst(20),
    I1 => cpi_d_inst(22),
    I2 => GRLFPC2_0_N_703_1,
    O => GRLFPC2_0_MOV_7_SQMUXA_3);
  x_grlfpc2_0_comb_fpdecode_mov5_1: LUT3 
  generic map(
    INIT => X"10"
  )
  port map (
    I0 => cpi_d_inst(9),
    I1 => cpi_d_inst(13),
    I2 => GRLFPC2_0_MOV_0_SQMUXA_2,
    O => GRLFPC2_0_COMB_FPDECODE_MOV5_1);
  x_grlfpc2_0_comb_fpdecode_un1_fpci_1_2: LUT4 
  generic map(
    INIT => X"0002"
  )
  port map (
    I0 => cpi_d_inst(5),
    I1 => cpi_d_inst(6),
    I2 => cpi_d_inst(9),
    I3 => cpi_d_inst(13),
    O => GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_1_0);
  x_grlfpc2_0_annulfpu_0_sqmuxa_1: LUT3 
  generic map(
    INIT => X"E0"
  )
  port map (
    I0 => cpi_e_annul,
    I1 => cpi_e_trap,
    I2 => GRLFPC2_0_R_E_FPOP,
    O => GRLFPC2_0_ANNULFPU_0_SQMUXA_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_sn_m3: LUT3 
  generic map(
    INIT => X"15"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_I(43),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_854);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_expybus_1_10x: LUT3 
  generic map(
    INIT => X"08"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(234),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_1(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_expybus_1_11x: LUT3 
  generic map(
    INIT => X"08"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(233),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_1(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_expybus_1_12x: LUT3 
  generic map(
    INIT => X"08"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(232),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_1(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_2_1x: LUT3 
  generic map(
    INIT => X"A8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_FAST(16),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(5),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzxbus_2_2x: LUT3 
  generic map(
    INIT => X"A8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_FAST(16),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(6),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sronemore: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(42),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(15),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un37_notxzyfromd: LUT4 
  generic map(
    INIT => X"0777"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(374),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(9),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(11),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(12),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTXZYFROMD_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_axb_12: LUT4 
  generic map(
    INIT => X"936C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1000,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_1(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_12);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_57: LUT4 
  generic map(
    INIT => X"8778"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(58),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(57),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_57);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_t_3_i_a2_0_0_0x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2281_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(375),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_T_3_I_A2_0_0(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathc_0_0: LUT3 
  generic map(
    INIT => X"01"
  )
  port map (
    I0 => GRLFPC2_0_R_MK_LDOP,
    I1 => GRLFPC2_0_R_MK_RST,
    I2 => GRLFPC2_0_R_MK_RST2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_2_0);
  x_grlfpc2_0_r_mk_ldopc_2: LUT3 
  generic map(
    INIT => X"01"
  )
  port map (
    I0 => cpi_d_annul,
    I1 => cpi_d_trap,
    I2 => cpi_flush,
    O => GRLFPC2_0_R_MK_LDOPC_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_entryshft_un9_s_11_1: LUT3 
  generic map(
    INIT => X"02"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(79),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(83),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(84),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN9_S_11_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_temp2: LUT3 
  generic map(
    INIT => X"10"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(65),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(71),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(75),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_r_dpath_inv_2: LUT4 
  generic map(
    INIT => X"0001"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(6),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_53_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_entryshft_un5_s_0: LUT3 
  generic map(
    INIT => X"01"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(78),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(84),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(85),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_aebeexc_un11_notbinfnan: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(247),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(248),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(249),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN11_NOTBINFNAN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_aebeexc_un11_notainfnan: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(234),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(235),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(236),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN11_NOTAINFNAN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_aebeexc_un5_notbzerodenorm: LUT3 
  generic map(
    INIT => X"01"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(247),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(248),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(249),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN5_NOTBZERODENORM_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_aebeexc_un5_notazerodenorm: LUT3 
  generic map(
    INIT => X"01"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(234),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(235),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(236),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN5_NOTAZERODENORM_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un5_xzybuslsbs: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(58),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(11),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN5_XZYBUSLSBS);
  x_grlfpc2_0_comb_un1_fpci: LUT3 
  generic map(
    INIT => X"01"
  )
  port map (
    I0 => cpi_flush,
    I1 => cpi_x_annul,
    I2 => cpi_x_trap,
    O => GRLFPC2_0_N_781);
  x_grlfpc2_0_comb_lockgen_un8_depcheck: LUT4_L 
  generic map(
    INIT => X"0001"
  )
  port map (
    I0 => GRLFPC2_0_R_A_LD,
    I1 => GRLFPC2_0_R_E_LD,
    I2 => GRLFPC2_0_R_M_LD,
    I3 => GRLFPC2_0_R_X_LD,
    LO => GRLFPC2_0_N_776);
  x_grlfpc2_0_comb_fpdecode_rs2d5_1: LUT3 
  generic map(
    INIT => X"04"
  )
  port map (
    I0 => cpi_d_inst(8),
    I1 => cpi_d_inst(9),
    I2 => cpi_d_inst(13),
    O => GRLFPC2_0_COMB_FPDECODE_RS2D5_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_feedbackmulxff_un18_feedback: LUT4 
  generic map(
    INIT => X"8000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(49),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(50),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(51),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(52),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN18_FEEDBACK);
  x_grlfpc2_0_comb_un1_fpci_3: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => cpi_a_cnt(1),
    I1 => GRLFPC2_0_R_A_RS1D,
    I2 => GRLFPC2_0_R_A_ST,
    O => GRLFPC2_0_COMB_UN1_FPCI_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_6_and_1: LUT3 
  generic map(
    INIT => X"01"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(50),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(52),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_6_AND_1);
  x_grlfpc2_0_comb_fpdecode_afq8_0: LUT4 
  generic map(
    INIT => X"0100"
  )
  port map (
    I0 => cpi_d_inst(20),
    I1 => cpi_d_inst(21),
    I2 => cpi_d_inst(22),
    I3 => cpi_d_inst(24),
    O => GRLFPC2_0_COMB_FPDECODE_AFQ8_0);
  x_grlfpc2_0_comb_fpdecode_un1_wren210_1_0_0: LUT3 
  generic map(
    INIT => X"20"
  )
  port map (
    I0 => cpi_d_inst(7),
    I1 => cpi_d_inst(8),
    I2 => cpi_d_inst(12),
    O => GRLFPC2_0_COMB_FPDECODE_UN1_WREN210_1_0_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_entryshft_s_cmp_0: LUT4 
  generic map(
    INIT => X"0040"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(79),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(82),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(84),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(85),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_S_CMP_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_entryshft_un14_s_mov_1: LUT3 
  generic map(
    INIT => X"02"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(80),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(81),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(82),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN14_S_MOV_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_wqstsets_1_4_6x: LUT4 
  generic map(
    INIT => X"0001"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(250),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(251),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(252),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(256),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_4(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_wqstsets_1_5_6x: LUT4 
  generic map(
    INIT => X"0001"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(253),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(254),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(255),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(257),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_5(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_wqstsets_1_4_5x: LUT4 
  generic map(
    INIT => X"0001"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(237),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(239),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(240),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(241),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_4(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_wqstsets_1_5_5x: LUT4 
  generic map(
    INIT => X"0001"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(238),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(242),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(243),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(244),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_5(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_aebeexc_un37_notainfnan_4: LUT4 
  generic map(
    INIT => X"8000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(237),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(238),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(239),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(240),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTAINFNAN_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_aebeexc_un37_notainfnan_5: LUT4 
  generic map(
    INIT => X"8000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(241),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(242),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(243),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(244),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTAINFNAN_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_aebeexc_un37_notbinfnan_4: LUT4 
  generic map(
    INIT => X"8000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(252),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(254),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(255),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(256),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTBINFNAN_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_aebeexc_un37_notbinfnan_5: LUT4 
  generic map(
    INIT => X"8000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(250),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(251),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(253),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(257),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTBINFNAN_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un21_notxzyfromd_i_0: LUT4_L 
  generic map(
    INIT => X"0777"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_DREG_FAST(53),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_FAST(375),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(11),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(13),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_I_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un4_notxzyfromd_i_0: LUT4 
  generic map(
    INIT => X"153F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_DREG_FAST(51),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_FAST(376),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(9),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(14),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_I_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_r_dpath_inv_6_1: LUT4 
  generic map(
    INIT => X"0001"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(7),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(9),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(10),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV_6_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un17_srtosticky_3: LUT4_L 
  generic map(
    INIT => X"0001"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(8),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(9),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN17_SRTOSTICKY_3);
  x_grlfpc2_0_r_mk_ldopc_1_0: LUT3 
  generic map(
    INIT => X"20"
  )
  port map (
    I0 => cpi_d_inst(23),
    I1 => cpi_d_inst(30),
    I2 => holdn,
    O => GRLFPC2_0_R_MK_LDOPC_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_52_trfwwbasiccell_un525_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(62),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_UN525_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_52_trfwwbasiccell_un354_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(62),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_UN354_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_52_trfwwbasiccell_un183_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(62),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_UN183_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_52_trfwwbasiccell_un12_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(62),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_UN12_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_49_trfwwbasiccell_un363_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(65),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_UN363_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_49_trfwwbasiccell_un534_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(65),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_UN534_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_36_trfwwbasiccell_un573_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(78),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_UN573_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_36_trfwwbasiccell_un402_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(78),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_UN402_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_36_trfwwbasiccell_un231_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(78),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_UN231_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_36_trfwwbasiccell_un60_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(78),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_UN60_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_15_trfwwbasiccell_un636_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(99),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_UN636_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_15_trfwwbasiccell_un465_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(99),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_UN465_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_15_trfwwbasiccell_un294_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(99),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_UN294_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_15_trfwwbasiccell_un123_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(99),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_UN123_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un2_mixoout3: LUT4 
  generic map(
    INIT => X"4450"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(7),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2008);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_Shift_3x: LUT2 
  generic map(
    INIT => X"6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_47_trfwwbasiccell_un540_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(67),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_UN540_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_47_trfwwbasiccell_un369_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(67),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_UN369_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_47_trfwwbasiccell_un198_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(67),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_UN198_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_14_trfwwbasiccell_un639_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(100),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_UN639_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_14_trfwwbasiccell_un468_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(100),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_UN468_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_14_trfwwbasiccell_un297_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(100),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_UN297_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_14_trfwwbasiccell_un126_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(100),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_UN126_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_13_trfwwbasiccell_un129_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(101),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_UN129_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_13_trfwwbasiccell_un300_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(101),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_UN300_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_13_trfwwbasiccell_un471_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(101),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_UN471_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_13_trfwwbasiccell_un642_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(101),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_UN642_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_0_trfwwbasiccell_un168_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(114),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_UN168_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_16_trfwwbasiccell_un633_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(98),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_UN633_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_19_trfwwbasiccell_un624_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(95),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_19_TRFWWBASICCELL_UN624_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_16_trfwwbasiccell_un462_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(98),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_UN462_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_16_trfwwbasiccell_un291_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(98),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_UN291_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_16_trfwwbasiccell_un120_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(98),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_UN120_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_19_trfwwbasiccell_un111_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(95),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_19_TRFWWBASICCELL_UN111_TEMP);
  x_grlfpc2_0_comb_dbgdata_5_29x: LUT4 
  generic map(
    INIT => X"3210"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => cpi_dbg_fsr,
    I2 => rfo1_data1(29),
    I3 => rfo2_data1(29),
    O => cpo_dbg_data(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_28_trfwwbasiccell_un597_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(86),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_UN597_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_28_trfwwbasiccell_un426_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(86),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_UN426_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_28_trfwwbasiccell_un255_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(86),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_UN255_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_28_trfwwbasiccell_un84_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(86),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_UN84_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_0_trfwwbasiccell_un510_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(114),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_UN510_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_0_trfwwbasiccell_un339_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(114),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_UN339_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_trfwwbasiccell_un651_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(104),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_UN651_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_trfwwbasiccell_un480_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(104),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_UN480_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_trfwwbasiccell_un309_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(104),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_UN309_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_trfwwbasiccell_un138_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(104),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_UN138_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_trfwwbasiccell_un648_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(103),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_UN648_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_trfwwbasiccell_un477_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(103),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_UN477_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_trfwwbasiccell_un306_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(103),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_UN306_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_trfwwbasiccell_un135_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(103),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_UN135_TEMP);
  x_grlfpc2_0_comb_dbgdata_5_28x: LUT4 
  generic map(
    INIT => X"3210"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => cpi_dbg_fsr,
    I2 => rfo1_data1(28),
    I3 => rfo2_data1(28),
    O => cpo_dbg_data(28));
  x_grlfpc2_0_comb_dbgdata_5_21x: LUT4 
  generic map(
    INIT => X"3210"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => cpi_dbg_fsr,
    I2 => rfo1_data1(21),
    I3 => rfo2_data1(21),
    O => cpo_dbg_data(21));
  x_grlfpc2_0_comb_dbgdata_5_20x: LUT4 
  generic map(
    INIT => X"3210"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => cpi_dbg_fsr,
    I2 => rfo1_data1(20),
    I3 => rfo2_data1(20),
    O => cpo_dbg_data(20));
  x_grlfpc2_0_comb_dbgdata_5_19x: LUT4 
  generic map(
    INIT => X"3210"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => cpi_dbg_fsr,
    I2 => rfo1_data1(19),
    I3 => rfo2_data1(19),
    O => cpo_dbg_data(19));
  x_grlfpc2_0_comb_dbgdata_5_15x: LUT4 
  generic map(
    INIT => X"3210"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => cpi_dbg_fsr,
    I2 => rfo1_data1(15),
    I3 => rfo2_data1(15),
    O => cpo_dbg_data(15));
  x_grlfpc2_0_comb_dbgdata_5_12x: LUT4 
  generic map(
    INIT => X"3210"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => cpi_dbg_fsr,
    I2 => rfo1_data1(12),
    I3 => rfo2_data1(12),
    O => cpo_dbg_data(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_Shift_1_0x: LUT4 
  generic map(
    INIT => X"99A5"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(25),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(57),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_Shift_2_1x: LUT4 
  generic map(
    INIT => X"99A5"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_Shift_3_2x: LUT4 
  generic map(
    INIT => X"99A5"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(5),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_trfwwbasiccell_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(58),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_55_trfwwbasiccell_un3_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(59),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_UN3_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_trfwwbasiccell_un6_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(60),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_UN6_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_53_trfwwbasiccell_un9_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(61),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_UN9_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_51_trfwwbasiccell_un15_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(63),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_UN15_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_50_trfwwbasiccell_un18_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_UN18_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_46_trfwwbasiccell_un30_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(68),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_UN30_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_45_trfwwbasiccell_un33_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(69),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_UN33_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_44_trfwwbasiccell_un36_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(70),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_UN36_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_43_trfwwbasiccell_un39_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(71),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_UN39_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_42_trfwwbasiccell_un42_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(72),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_UN42_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_41_trfwwbasiccell_un45_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(73),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_UN45_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_40_trfwwbasiccell_un48_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(74),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_UN48_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_39_trfwwbasiccell_un51_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_UN51_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_38_trfwwbasiccell_un54_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_UN54_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_37_trfwwbasiccell_un57_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(77),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_UN57_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_35_trfwwbasiccell_un63_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(79),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_UN63_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_34_trfwwbasiccell_un66_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(80),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_UN66_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_33_trfwwbasiccell_un69_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(81),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_UN69_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_32_trfwwbasiccell_un72_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(82),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_UN72_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_31_trfwwbasiccell_un75_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_UN75_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_30_trfwwbasiccell_un78_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(84),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_UN78_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_29_trfwwbasiccell_un81_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(85),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_UN81_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_27_trfwwbasiccell_un87_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(87),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_UN87_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_26_trfwwbasiccell_un90_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(88),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_UN90_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_25_trfwwbasiccell_un93_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(89),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_UN93_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_trfwwbasiccell_un96_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(90),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_UN96_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_trfwwbasiccell_un99_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(91),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_UN99_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_22_trfwwbasiccell_un102_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(92),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_UN102_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_21_trfwwbasiccell_un105_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(93),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_UN105_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_20_trfwwbasiccell_un108_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(94),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_UN108_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_18_trfwwbasiccell_un114_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(96),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_18_TRFWWBASICCELL_UN114_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_17_trfwwbasiccell_un117_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(97),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_UN117_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_12_trfwwbasiccell_un132_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(102),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_UN132_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_trfwwbasiccell_un141_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(105),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_UN141_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_8_trfwwbasiccell_un144_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(106),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_UN144_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_trfwwbasiccell_un147_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(107),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_UN147_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_6_trfwwbasiccell_un150_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(108),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_UN150_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_5_trfwwbasiccell_un153_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(109),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_UN153_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_trfwwbasiccell_un156_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(110),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_UN156_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_trfwwbasiccell_un159_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(111),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_UN159_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_trfwwbasiccell_un162_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(112),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_UN162_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_1_trfwwbasiccell_un165_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(113),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_UN165_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_trfwwbasiccell_un171_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(58),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_UN171_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_55_trfwwbasiccell_un174_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(59),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_UN174_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_trfwwbasiccell_un177_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(60),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_UN177_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_53_trfwwbasiccell_un180_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(61),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_UN180_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_51_trfwwbasiccell_un186_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(63),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_UN186_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_46_trfwwbasiccell_un201_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(68),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_UN201_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_45_trfwwbasiccell_un204_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(69),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_UN204_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_44_trfwwbasiccell_un207_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(70),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_UN207_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_43_trfwwbasiccell_un210_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(71),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_UN210_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_41_trfwwbasiccell_un216_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(73),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_UN216_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_40_trfwwbasiccell_un219_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(74),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_UN219_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_39_trfwwbasiccell_un222_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_UN222_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_38_trfwwbasiccell_un225_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_UN225_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_37_trfwwbasiccell_un228_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(77),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_UN228_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_35_trfwwbasiccell_un234_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(79),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_UN234_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_34_trfwwbasiccell_un237_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(80),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_UN237_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_33_trfwwbasiccell_un240_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(81),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_UN240_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_32_trfwwbasiccell_un243_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(82),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_UN243_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_31_trfwwbasiccell_un246_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_UN246_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_29_trfwwbasiccell_un252_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(85),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_UN252_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_27_trfwwbasiccell_un258_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(87),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_UN258_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_26_trfwwbasiccell_un261_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(88),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_UN261_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_25_trfwwbasiccell_un264_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(89),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_UN264_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_trfwwbasiccell_un267_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(90),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_UN267_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_trfwwbasiccell_un270_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(91),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_UN270_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_22_trfwwbasiccell_un273_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(92),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_UN273_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_21_trfwwbasiccell_un276_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(93),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_UN276_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_17_trfwwbasiccell_un288_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(97),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_UN288_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_12_trfwwbasiccell_un303_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(102),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_UN303_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_trfwwbasiccell_un312_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(105),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_UN312_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_8_trfwwbasiccell_un315_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(106),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_UN315_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_trfwwbasiccell_un318_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(107),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_UN318_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_6_trfwwbasiccell_un321_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(108),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_UN321_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_5_trfwwbasiccell_un324_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(109),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_UN324_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_trfwwbasiccell_un327_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(110),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_UN327_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_trfwwbasiccell_un330_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(111),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_UN330_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_trfwwbasiccell_un333_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(112),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_UN333_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_1_trfwwbasiccell_un336_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(113),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_UN336_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_trfwwbasiccell_un342_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(58),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_UN342_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_55_trfwwbasiccell_un345_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(59),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_UN345_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_trfwwbasiccell_un348_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(60),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_UN348_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_53_trfwwbasiccell_un351_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(61),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_UN351_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_51_trfwwbasiccell_un357_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(63),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_UN357_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_50_trfwwbasiccell_un360_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_UN360_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_48_trfwwbasiccell_un366_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_UN366_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_46_trfwwbasiccell_un372_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(68),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_UN372_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_45_trfwwbasiccell_un375_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(69),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_UN375_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_44_trfwwbasiccell_un378_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(70),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_UN378_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_43_trfwwbasiccell_un381_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(71),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_UN381_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_42_trfwwbasiccell_un384_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(72),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_UN384_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_41_trfwwbasiccell_un387_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(73),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_UN387_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_40_trfwwbasiccell_un390_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(74),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_UN390_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_39_trfwwbasiccell_un393_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_UN393_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_38_trfwwbasiccell_un396_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_UN396_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_37_trfwwbasiccell_un399_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(77),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_UN399_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_35_trfwwbasiccell_un405_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(79),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_UN405_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_34_trfwwbasiccell_un408_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(80),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_UN408_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_33_trfwwbasiccell_un411_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(81),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_UN411_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_32_trfwwbasiccell_un414_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(82),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_UN414_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_31_trfwwbasiccell_un417_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_UN417_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_30_trfwwbasiccell_un420_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(84),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_UN420_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_29_trfwwbasiccell_un423_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(85),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_UN423_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_27_trfwwbasiccell_un429_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(87),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_UN429_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_26_trfwwbasiccell_un432_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(88),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_UN432_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_25_trfwwbasiccell_un435_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(89),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_UN435_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_trfwwbasiccell_un438_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(90),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_UN438_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_trfwwbasiccell_un441_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(91),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_UN441_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_22_trfwwbasiccell_un444_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(92),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_UN444_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_21_trfwwbasiccell_un447_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(93),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_UN447_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_20_trfwwbasiccell_un450_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(94),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_UN450_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_17_trfwwbasiccell_un459_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(97),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_UN459_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_12_trfwwbasiccell_un474_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(102),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_UN474_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_trfwwbasiccell_un483_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(105),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_UN483_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_8_trfwwbasiccell_un486_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(106),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_UN486_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_trfwwbasiccell_un489_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(107),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_UN489_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_6_trfwwbasiccell_un492_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(108),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_UN492_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_5_trfwwbasiccell_un495_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(109),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_UN495_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_trfwwbasiccell_un498_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(110),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_UN498_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_trfwwbasiccell_un501_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(111),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_UN501_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_trfwwbasiccell_un504_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(112),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_UN504_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_1_trfwwbasiccell_un507_temp: LUT4 
  generic map(
    INIT => X"5A3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(113),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_UN507_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_trfwwbasiccell_un513_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(58),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_UN513_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_55_trfwwbasiccell_un516_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(59),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_UN516_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_trfwwbasiccell_un519_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(60),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_UN519_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_53_trfwwbasiccell_un522_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(61),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_UN522_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_51_trfwwbasiccell_un528_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(63),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_UN528_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_50_trfwwbasiccell_un531_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_UN531_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_48_trfwwbasiccell_un537_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_UN537_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_46_trfwwbasiccell_un543_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(68),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_UN543_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_45_trfwwbasiccell_un546_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(69),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_UN546_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_44_trfwwbasiccell_un549_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(70),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_UN549_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_43_trfwwbasiccell_un552_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(71),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_UN552_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_42_trfwwbasiccell_un555_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(72),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_UN555_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_41_trfwwbasiccell_un558_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(73),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_UN558_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_40_trfwwbasiccell_un561_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(74),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_UN561_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_37_trfwwbasiccell_un570_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(77),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_UN570_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_35_trfwwbasiccell_un576_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(79),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_UN576_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_34_trfwwbasiccell_un579_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(80),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_UN579_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_33_trfwwbasiccell_un582_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(81),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_UN582_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_32_trfwwbasiccell_un585_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(82),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_UN585_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_31_trfwwbasiccell_un588_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_UN588_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_30_trfwwbasiccell_un591_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(84),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_UN591_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_29_trfwwbasiccell_un594_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(85),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_UN594_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_27_trfwwbasiccell_un600_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(87),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_UN600_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_26_trfwwbasiccell_un603_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(88),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_UN603_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_25_trfwwbasiccell_un606_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(89),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_UN606_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_trfwwbasiccell_un609_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(90),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_UN609_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_trfwwbasiccell_un612_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(91),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_UN612_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_22_trfwwbasiccell_un615_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(92),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_UN615_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_21_trfwwbasiccell_un618_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(93),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_UN618_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_20_trfwwbasiccell_un621_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(94),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_UN621_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_18_trfwwbasiccell_un627_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(96),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_18_TRFWWBASICCELL_UN627_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_17_trfwwbasiccell_un630_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(97),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_UN630_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_12_trfwwbasiccell_un645_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(102),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_UN645_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_trfwwbasiccell_un654_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(105),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_UN654_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_8_trfwwbasiccell_un657_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(106),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_UN657_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_trfwwbasiccell_un660_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(107),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_UN660_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_6_trfwwbasiccell_un663_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(108),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_UN663_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_5_trfwwbasiccell_un666_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(109),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_UN666_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_trfwwbasiccell_un669_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(110),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_UN669_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_trfwwbasiccell_un672_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(111),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_UN672_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_trfwwbasiccell_un675_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(112),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_UN675_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_1_trfwwbasiccell_un678_temp: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(113),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_UN678_TEMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_expybus_1_4x: LUT4 
  generic map(
    INIT => X"C0A0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(240),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_1(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_3x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(112),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_16_REP1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_FAST(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_4x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(111),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_16_REP1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_FAST(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_5x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(110),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_16_REP1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_FAST(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_6x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(109),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_16_REP1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_FAST(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_7x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(108),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_16_REP1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_FAST(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_8x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(107),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_16_REP1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_FAST(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_9x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(106),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_16_REP1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_FAST(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_10x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(105),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_16_REP1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_FAST(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_13x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(102),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_FAST(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_18x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(97),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_19x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(96),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_21x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(94),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_22x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(93),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_23x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(92),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_24x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(91),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_25x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(90),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_26x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(89),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_27x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(88),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_28x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(87),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_30x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(85),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_31x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(84),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_0_0x: LUT3 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(15),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_0_1x: LUT3 
  generic map(
    INIT => X"8C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(15),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_0_2x: LUT3 
  generic map(
    INIT => X"8C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(15),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srcontrol_1_0_3x: LUT4 
  generic map(
    INIT => X"8BCF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_I(43),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(15),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_ss6_0: LUT3 
  generic map(
    INIT => X"BA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(7),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(9),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SS6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_1_0_2x: LUT4 
  generic map(
    INIT => X"FCAA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(242),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(30),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_846);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_expybus_1_0_0_5x: LUT4 
  generic map(
    INIT => X"C0AA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(239),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(30),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1017);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_12x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(103),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_16_REP1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_FAST(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_11x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(104),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_16_REP1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_FAST(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_29x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(86),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_20x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(95),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_17x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(98),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_FAST(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_14x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(101),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_FAST(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_15x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(100),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_FAST(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_16x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(99),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_FAST(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_57: LUT4 
  generic map(
    INIT => X"E4D7"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(58),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_I(19),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_57);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_42_0: LUT3 
  generic map(
    INIT => X"87"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(73),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_42_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_44_0: LUT3 
  generic map(
    INIT => X"87"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(71),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_44_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_waitq_i_0x: LUT3 
  generic map(
    INIT => X"47"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(58),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_I(19),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I(0));
  x_grlfpc2_0_v_state_1_sqmuxa_1: LUT3 
  generic map(
    INIT => X"13"
  )
  port map (
    I0 => GRLFPC2_0_R_X_AFQ,
    I1 => GRLFPC2_0_R_X_SEQERR,
    I2 => GRLFPC2_0_SEQERR_1_SQMUXA_1_SN,
    O => GRLFPC2_0_V_STATE_1_SQMUXA_1);
  x_grlfpc2_0_v_fsr_ftt_1_sqmuxa_2_2: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_N_781,
    I1 => GRLFPC2_0_R_X_SEQERR,
    O => GRLFPC2_0_V_FSR_FTT_1_SQMUXA_2_2);
  x_grlfpc2_0_wren2_1_sqmuxa_1: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_N_781,
    I1 => GRLFPC2_0_R_X_SEQERR,
    O => GRLFPC2_0_WREN2_1_SQMUXA_1);
  x_grlfpc2_0_v_i_exec_0_sqmuxa: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_N_781,
    I1 => GRLFPC2_0_R_X_FPOP,
    O => GRLFPC2_0_V_I_EXEC_0_SQMUXA);
  x_grlfpc2_0_wraddr_0_sqmuxa_1: LUT3 
  generic map(
    INIT => X"20"
  )
  port map (
    I0 => GRLFPC2_0_N_781,
    I1 => GRLFPC2_0_R_X_AFSR,
    I2 => GRLFPC2_0_R_X_LD,
    O => GRLFPC2_0_WRADDR_0_SQMUXA_1);
  x_grlfpc2_0_comb_fpdecode_un3_op: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => cpi_d_inst(23),
    I1 => GRLFPC2_0_MOV_7_SQMUXA_3,
    O => GRLFPC2_0_COMB_FPDECODE_UN3_OP);
  x_grlfpc2_0_comb_fpdecode_afq3: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => cpi_d_inst(19),
    I1 => cpi_d_inst(20),
    I2 => GRLFPC2_0_COMB_FPDECODE_AFQ4_1,
    O => GRLFPC2_0_COMB_FPDECODE_AFQ3);
  x_grlfpc2_0_comb_un1_r_a_rs1_1: LUT3 
  generic map(
    INIT => X"51"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN1_FPCI_3,
    I1 => GRLFPC2_0_R_A_RS1(0),
    I2 => GRLFPC2_0_R_A_RS1D,
    O => GRLFPC2_0_N_772);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_condmuxmulxff_un4_notsqrtlftcc: LUT4 
  generic map(
    INIT => X"0054"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(65),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(75),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(76),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(77),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CONDMUXMULXFF_UN4_NOTSQRTLFTCC);
  x_grlfpc2_0_comb_fpdecode_afq7: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => cpi_d_inst(19),
    I1 => cpi_d_inst(20),
    I2 => GRLFPC2_0_COMB_FPDECODE_AFQ7_1,
    O => GRLFPC2_0_COMB_FPDECODE_AFQ7);
  x_grlfpc2_0_v_fsr_nonstd_0_sqmuxa_2: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_N_781,
    I1 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA,
    O => GRLFPC2_0_V_FSR_AEXC_1_SQMUXA_SN);
  x_grlfpc2_0_comb_un1_fpci_4: LUT3 
  generic map(
    INIT => X"51"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN1_FPCI_3,
    I1 => GRLFPC2_0_R_A_RS2(0),
    I2 => GRLFPC2_0_R_A_RS2D,
    O => GRLFPC2_0_N_771);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un46_xzybuslsbs: LUT2 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTXZYFROMD_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(231),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN46_XZYBUSLSBS);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un3_inexact: LUT3 
  generic map(
    INIT => X"2A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_NOTAM2_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(54),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN3_INEXACT);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_mixoIn_3_0_1x: LUT3 
  generic map(
    INIT => X"5C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(372),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un4_temp_2_0_am_0x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(54),
    LO => N_12084);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_4x: LUT4 
  generic map(
    INIT => X"ACA0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_992,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(4));
  x_grlfpc2_0_comb_dbgdata_5_0_0x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_fsr,
    I1 => GRLFPC2_0_N_311,
    I2 => GRLFPC2_0_R_FSR_CEXC(0),
    O => cpo_dbg_data(0));
  x_grlfpc2_0_comb_dbgdata_5_0_1x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_fsr,
    I1 => GRLFPC2_0_N_312,
    I2 => GRLFPC2_0_R_FSR_CEXC(1),
    O => cpo_dbg_data(1));
  x_grlfpc2_0_comb_dbgdata_5_0_2x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_fsr,
    I1 => GRLFPC2_0_N_313,
    I2 => GRLFPC2_0_R_FSR_CEXC(2),
    O => cpo_dbg_data(2));
  x_grlfpc2_0_comb_dbgdata_5_0_3x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_fsr,
    I1 => GRLFPC2_0_N_314,
    I2 => GRLFPC2_0_R_FSR_CEXC(3),
    O => cpo_dbg_data(3));
  x_grlfpc2_0_comb_dbgdata_5_0_5x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_fsr,
    I1 => GRLFPC2_0_N_316,
    I2 => GRLFPC2_0_R_FSR_AEXC(0),
    O => cpo_dbg_data(5));
  x_grlfpc2_0_comb_dbgdata_5_0_6x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_fsr,
    I1 => GRLFPC2_0_N_317,
    I2 => GRLFPC2_0_R_FSR_AEXC(1),
    O => cpo_dbg_data(6));
  x_grlfpc2_0_comb_dbgdata_5_0_7x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_fsr,
    I1 => GRLFPC2_0_N_318,
    I2 => GRLFPC2_0_R_FSR_AEXC(2),
    O => cpo_dbg_data(7));
  x_grlfpc2_0_comb_dbgdata_5_0_8x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_fsr,
    I1 => GRLFPC2_0_N_319,
    I2 => GRLFPC2_0_R_FSR_AEXC(3),
    O => cpo_dbg_data(8));
  x_grlfpc2_0_comb_dbgdata_5_0_9x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_fsr,
    I1 => GRLFPC2_0_N_320,
    I2 => GRLFPC2_0_R_FSR_AEXC(4),
    O => cpo_dbg_data(9));
  x_grlfpc2_0_comb_dbgdata_5_0_10x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => cpi_dbg_fsr,
    I1 => CPO_CC_0_INT_3,
    I2 => GRLFPC2_0_N_321,
    O => cpo_dbg_data(10));
  x_grlfpc2_0_comb_dbgdata_5_0_11x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => cpi_dbg_fsr,
    I1 => CPO_CC_1_INT_4,
    I2 => GRLFPC2_0_N_322,
    O => cpo_dbg_data(11));
  x_grlfpc2_0_comb_dbgdata_5_0_22x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_fsr,
    I1 => GRLFPC2_0_N_333,
    I2 => GRLFPC2_0_R_FSR_NONSTD,
    O => cpo_dbg_data(22));
  x_grlfpc2_0_comb_dbgdata_5_0_23x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_fsr,
    I1 => GRLFPC2_0_N_334,
    I2 => GRLFPC2_0_R_FSR_TEM(0),
    O => cpo_dbg_data(23));
  x_grlfpc2_0_comb_dbgdata_5_0_24x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_fsr,
    I1 => GRLFPC2_0_N_335,
    I2 => GRLFPC2_0_R_FSR_TEM(1),
    O => cpo_dbg_data(24));
  x_grlfpc2_0_comb_dbgdata_5_0_25x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_fsr,
    I1 => GRLFPC2_0_N_336,
    I2 => GRLFPC2_0_R_FSR_TEM(2),
    O => cpo_dbg_data(25));
  x_grlfpc2_0_comb_dbgdata_5_0_27x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_fsr,
    I1 => GRLFPC2_0_N_338,
    I2 => GRLFPC2_0_R_FSR_TEM(4),
    O => cpo_dbg_data(27));
  x_grlfpc2_0_comb_dbgdata_5_0_30x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_fsr,
    I1 => GRLFPC2_0_N_341,
    I2 => GRLFPC2_0_R_FSR_RD(0),
    O => cpo_dbg_data(30));
  x_grlfpc2_0_comb_dbgdata_5_0_31x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_fsr,
    I1 => GRLFPC2_0_N_342,
    I2 => GRLFPC2_0_R_FSR_RD(1),
    O => cpo_dbg_data(31));
  x_grlfpc2_0_comb_dbgdata_5_1_14x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_fsr,
    I1 => GRLFPC2_0_N_325,
    I2 => GRLFPC2_0_R_FSR_FTT(0),
    O => cpo_dbg_data(14));
  x_grlfpc2_0_comb_dbgdata_5_1_4x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_fsr,
    I1 => GRLFPC2_0_N_315,
    I2 => GRLFPC2_0_R_FSR_CEXC(4),
    O => cpo_dbg_data(4));
  x_grlfpc2_0_comb_dbgdata_5_1_am_13x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => rfo1_data1(13),
    I2 => rfo2_data1(13),
    O => N_12086);
  x_grlfpc2_0_comb_dbgdata_5_1_bm_13x: LUT2 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => GRLFPC2_0_R_STATE(0),
    I1 => GRLFPC2_0_R_STATE(1),
    O => N_12087);
  x_grlfpc2_0_comb_dbgdata_5_1_13x: MUXF5 port map (
      I0 => N_12086,
      I1 => N_12087,
      S => cpi_dbg_fsr,
      O => cpo_dbg_data(13));
  x_grlfpc2_0_comb_dbgdata_5_1_26x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_fsr,
    I1 => GRLFPC2_0_N_337,
    I2 => GRLFPC2_0_R_FSR_TEM(3),
    O => cpo_dbg_data(26));
  x_grlfpc2_0_comb_dbgdata_5_1_16x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_dbg_fsr,
    I1 => GRLFPC2_0_N_327,
    I2 => GRLFPC2_0_R_FSR_FTT(2),
    O => cpo_dbg_data(16));
  x_grlfpc2_0_annulres_0_sqmuxa_3_0: LUT4_L 
  generic map(
    INIT => X"E000"
  )
  port map (
    I0 => cpi_a_annul,
    I1 => cpi_a_trap,
    I2 => GRLFPC2_0_ANNULRES_0_SQMUXA_3_2,
    I3 => GRLFPC2_0_R_A_FPOP,
    LO => GRLFPC2_0_ANNULRES_0_SQMUXA_3_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un1_mifrominst_0: LUT3 
  generic map(
    INIT => X"02"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(63),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(77),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN1_MIFROMINST_0);
  x_grlfpc2_0_fpi_ldop: LUT4 
  generic map(
    INIT => X"0100"
  )
  port map (
    I0 => GRLFPC2_0_R_MK_LDOP,
    I1 => GRLFPC2_0_R_MK_RST,
    I2 => GRLFPC2_0_R_MK_RST2,
    I3 => rst,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0);
  x_grlfpc2_0_I_251: LUT4 
  generic map(
    INIT => X"1000"
  )
  port map (
    I0 => cpi_a_annul,
    I1 => cpi_a_trap,
    I2 => GRLFPC2_0_R_A_FPOP,
    I3 => GRLFPC2_0_R_A_MOV,
    O => GRLFPC2_0_N_691);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_entryshft_s_cmp: LUT3_L 
  generic map(
    INIT => X"08"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_S_CMP_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_ENTRYSHFT_S_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(78),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_S_CMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un15_wqstsets: LUT4 
  generic map(
    INIT => X"1000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(4),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(42),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(15),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1991);
  x_grlfpc2_0_comb_lockgen_depcheck: LUT4 
  generic map(
    INIT => X"0002"
  )
  port map (
    I0 => GRLFPC2_0_ANNULRES_0_SQMUXA_3_2,
    I1 => GRLFPC2_0_R_A_FPOP,
    I2 => GRLFPC2_0_R_I_EXEC,
    I3 => GRLFPC2_0_R_X_FPOP,
    O => GRLFPC2_0_N_777);
  x_grlfpc2_0_mov_2_sqmuxa_1_1: LUT4 
  generic map(
    INIT => X"0400"
  )
  port map (
    I0 => cpi_d_inst(9),
    I1 => cpi_d_inst(10),
    I2 => cpi_d_inst(13),
    I3 => GRLFPC2_0_MOV_0_SQMUXA_3,
    O => GRLFPC2_0_MOV_2_SQMUXA_1_1);
  x_grlfpc2_0_comb_un8_ccv_1: LUT4 
  generic map(
    INIT => X"0013"
  )
  port map (
    I0 => cpi_e_inst(19),
    I1 => GRLFPC2_0_COMB_UN22_CCV,
    I2 => GRLFPC2_0_R_E_FPOP,
    I3 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA,
    O => GRLFPC2_0_COMB_UN8_CCV_1);
  x_grlfpc2_0_comb_lock_1_1_0: LUT4 
  generic map(
    INIT => X"0001"
  )
  port map (
    I0 => cpi_d_annul,
    I1 => cpi_d_trap,
    I2 => GRLFPC2_0_R_STATE(0),
    I3 => GRLFPC2_0_R_STATE(1),
    O => GRLFPC2_0_COMB_LOCK_1_1_0);
  x_grlfpc2_0_comb_annulfpu_1_u_0: LUT4_L 
  generic map(
    INIT => X"010F"
  )
  port map (
    I0 => cpi_a_annul,
    I1 => cpi_a_trap,
    I2 => GRLFPC2_0_ANNULFPU_0_SQMUXA_1,
    I3 => GRLFPC2_0_R_A_FPOP,
    LO => GRLFPC2_0_COMB_ANNULFPU_1_U_0);
  x_grlfpc2_0_comb_un1_mexc_2: LUT3 
  generic map(
    INIT => X"01"
  )
  port map (
    I0 => GRLFPC2_0_COMB_MEXC_1(2),
    I1 => GRLFPC2_0_COMB_MEXC_1(3),
    I2 => GRLFPC2_0_COMB_MEXC_1(4),
    O => GRLFPC2_0_COMB_UN1_MEXC_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_entryshft_un4_s_sqrt_1_0: LUT4 
  generic map(
    INIT => X"0200"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_ENTRYSHFT_S_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(78),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(82),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(85),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN4_S_SQRT_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_53x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(62),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(262),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_57x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(58),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(258),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_16x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(99),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(299),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_48x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(67),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(267),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_14x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(101),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(301),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_2x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(113),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(313),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_3x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(112),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(312),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_5x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(110),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(310),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_6x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(109),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(309),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_20x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(95),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(295),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_22x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(93),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(293),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_17x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(98),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(298),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_52x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(63),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(263),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_15x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(100),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(300),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_44x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(71),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(271),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m2_0x: LUT3 
  generic map(
    INIT => X"BA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(15),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M2(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_29x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(86),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(286),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_temp_2_0x: LUT3 
  generic map(
    INIT => X"0E"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_2(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_54x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(61),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(261),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_56x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(59),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(259),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_37x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(78),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(278),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_39x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(276),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_40x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(275),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_46x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(69),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(269),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_47x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(68),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(268),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_19x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(96),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(296),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_21x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(94),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(294),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_9x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(106),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(306),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_12x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(103),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(303),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_26x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(89),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(289),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_32x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(283),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_18x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(97),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(297),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_expybus_1_6x: LUT4 
  generic map(
    INIT => X"A0C0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPYBUS_2(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(238),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_1(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_55x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(60),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(260),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_51x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(264),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_50x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(65),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(265),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_49x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(266),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_45x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(70),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(270),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_43x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(72),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(272),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_42x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(73),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(273),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_41x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(74),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(274),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_38x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(77),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(277),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_36x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(79),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(279),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_35x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(80),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(280),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_34x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(81),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(281),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_33x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(82),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(282),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_31x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(84),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(284),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_30x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(85),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(285),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_28x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(87),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(287),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_27x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(88),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(288),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_25x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(90),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(290),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_24x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(91),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(291),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_23x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(92),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(292),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_13x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(102),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(302),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_11x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(104),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(304),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_10x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(105),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(305),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_8x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(107),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(307),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_7x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(108),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(308),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_4x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(111),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(311),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlxershft_SumIn_4_1x: LUT4 
  generic map(
    INIT => X"11F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(114),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(314),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_113x: LUT2 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2008,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(113));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_temp_1_0x: LUT3 
  generic map(
    INIT => X"0E"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_2x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(113),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_FAST(17),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_1_0_1x: LUT3 
  generic map(
    INIT => X"5C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2016,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(243),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_845);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_1_0_3x: LUT3 
  generic map(
    INIT => X"5C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2017,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(241),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_847);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_am_2x: LUT3 
  generic map(
    INIT => X"E0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
    O => N_12088);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_bm_2x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(242),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(255),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
    O => N_12089);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_2x: MUXF5 port map (
      I0 => N_12088,
      I1 => N_12089,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_am_5x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
    O => N_12090);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_bm_5x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(239),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(252),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
    O => N_12091);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_5x: MUXF5 port map (
      I0 => N_12090,
      I1 => N_12091,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_am_6x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
    O => N_12092);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_bm_6x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(238),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(251),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
    O => N_12093);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_6x: MUXF5 port map (
      I0 => N_12092,
      I1 => N_12093,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_expybus_1_0_0_7x: LUT4 
  generic map(
    INIT => X"0CAC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPYBUS_2(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(237),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1019);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_expybus_1_0_0_8x: LUT4 
  generic map(
    INIT => X"0CAC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPYBUS_2(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(236),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1020);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_expybus_1_0_0_9x: LUT4 
  generic map(
    INIT => X"0CAC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPYBUS_2(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(235),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1021);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_1x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(114),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_FAST(17),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(1));
  x_grlfpc2_0_comb_isfpop2_1_0: LUT3 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => cpi_x_inst(19),
    I1 => GRLFPC2_0_COMB_UN1_R_I_V,
    I2 => GRLFPC2_0_R_I_INST(19),
    O => GRLFPC2_0_COMB_ISFPOP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_1_0_0x: LUT3 
  generic map(
    INIT => X"5C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_COMPUTECONST_UN49_RESVEC,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(244),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_844);
  x_grlfpc2_0_comb_annulfpu_1_0_0: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_N_781,
    I1 => GRLFPC2_0_R_X_FPOP,
    I2 => GRLFPC2_0_R_X_SEQERR,
    O => GRLFPC2_0_N_206);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzxbus_0_0x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(115),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_FAST(17),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_16_0: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(99),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_16_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_23_0: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(92),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_23_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_19_0: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(96),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_19_0);
  x_grlfpc2_0_comb_N_712_i: LUT4 
  generic map(
    INIT => X"FEDC"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => cpi_dbg_fsr,
    I2 => rfo1_data1(17),
    I3 => rfo2_data1(17),
    O => cpo_dbg_data(17));
  x_grlfpc2_0_comb_N_711_i: LUT4 
  generic map(
    INIT => X"FEDC"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => cpi_dbg_fsr,
    I2 => rfo1_data1(18),
    I3 => rfo2_data1(18),
    O => cpo_dbg_data(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un39_xzybuslsbs: LUT4 
  generic map(
    INIT => X"7050"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(57),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(10),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN39_XZYBUSLSBS);
  x_grlfpc2_0_comb_v_a_afsr_1_m0_0: LUT4 
  generic map(
    INIT => X"8CAF"
  )
  port map (
    I0 => cpi_d_inst(20),
    I1 => cpi_d_inst(23),
    I2 => GRLFPC2_0_COMB_FPDECODE_AFQ4_1,
    I3 => GRLFPC2_0_COMB_FPDECODE_AFQ8_0,
    O => GRLFPC2_0_N_716);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_un1_u_snnotdb: LUT2 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN1_U_SNNOTDB);
  x_grlfpc2_0_v_state_1_sqmuxa: LUT3 
  generic map(
    INIT => X"70"
  )
  port map (
    I0 => cpi_dbg_data(28),
    I1 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
    I2 => rst,
    O => GRLFPC2_0_V_STATE_1_SQMUXA);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_un12_u_snnotdb_1: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(65),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN12_U_SNNOTDB_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_m_1_51x: LUT2 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_srtosticky_1: LUT4 
  generic map(
    INIT => X"FD00"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN17_SRTOSTICKY_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(10),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(11),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlbregexp_ExpBregLC_1_1x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(25),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_EXPBREGLC_1(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_SignResult: LUT4 
  generic map(
    INIT => X"B51F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2031,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_AREGXORBREG,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(23),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(12),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2000);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_29_trfwwbasiccell_temp2_1_0: LUT4 
  generic map(
    INIT => X"D872"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_UN252_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(84),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_30_trfwwbasiccell_temp2_1_0: LUT4 
  generic map(
    INIT => X"C693"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(84),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_41_trfwwbasiccell_temp2_2_0: LUT4 
  generic map(
    INIT => X"D872"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_UN216_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(72),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_39_trfwwbasiccell_temp2_2_0: LUT4 
  generic map(
    INIT => X"C693"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(74),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_47_trfwwbasiccell_temp2_1_0: LUT4_L 
  generic map(
    INIT => X"C693"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(67),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_46_trfwwbasiccell_temp2_0: LUT4_L 
  generic map(
    INIT => X"D872"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_UN30_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(67),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_18_trfwwbasiccell_temp2_0: LUT4 
  generic map(
    INIT => X"C693"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(95),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(96),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_18_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_42_trfwwbasiccell_temp2_2_0: LUT4 
  generic map(
    INIT => X"C693"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(71),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(72),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_37_trfwwbasiccell_temp2_1_0: LUT4 
  generic map(
    INIT => X"D872"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_UN570_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_38_trfwwbasiccell_temp2_2_0: LUT4 
  generic map(
    INIT => X"C693"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_18_trfwwbasiccell_temp2_2_0: LUT4 
  generic map(
    INIT => X"C693"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(95),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(96),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_18_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_48_trfwwbasiccell_temp2_2_0: LUT4_L 
  generic map(
    INIT => X"C693"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(65),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_TEMP2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_trfwwbasiccell_temp2_3_0: LUT3 
  generic map(
    INIT => X"63"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(58),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_19_trfwwbasiccell_temp2_3_0: LUT4 
  generic map(
    INIT => X"C693"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(94),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(95),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_19_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_1x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(48),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_2x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(47),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_3x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(46),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(54),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_4x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(45),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_5x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(44),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(52),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_6x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(43),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_7x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(50),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_10x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(47),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_11x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(38),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(46),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_12x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(37),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(45),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_13x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(36),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(44),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_14x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(35),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(43),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_15x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(34),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(42),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_18x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(31),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(39),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_19x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(38),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_20x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(37),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_21x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(28),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_22x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(27),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(35),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_23x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(26),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(34),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_24x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(25),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(33),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_25x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(24),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(32),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_26x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(31),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_27x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(22),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(30),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_28x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(29),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_30x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(27),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_31x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(18),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(26),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_32x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(25),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_33x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(24),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_34x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(15),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_35x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(14),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(22),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_39x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(10),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(18),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_40x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(9),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_42x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(15),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_43x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(14),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_44x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(13),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_47x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(10),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_48x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(9),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_50x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(3),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_51x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_52x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(5),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_54x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_55x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(8),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_56x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(8),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_57x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(8),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_41x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(16),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_49x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_20_trfwwbasiccell_temp2_1_0: LUT4 
  generic map(
    INIT => X"C693"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(93),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(94),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_49_trfwwbasiccell_temp2_0: LUT4_L 
  generic map(
    INIT => X"C693"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(65),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_15_trfwwbasiccell_temp2_3_0: LUT4_L 
  generic map(
    INIT => X"F690"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(4),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_UN465_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_UN462_TEMP,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_17_trfwwbasiccell_temp2_0: LUT4 
  generic map(
    INIT => X"D872"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_UN288_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(96),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_47_trfwwbasiccell_temp2_0: LUT4 
  generic map(
    INIT => X"D872"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_UN198_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_0_trfwwbasiccell_temp2_3_0: LUT4 
  generic map(
    INIT => X"C693"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(113),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(114),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_0x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(49),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(57),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_9x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(48),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_8x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(41),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(49),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_17_trfwwbasiccell_temp2_3_0: LUT4 
  generic map(
    INIT => X"D872"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_UN459_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(96),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_TEMP2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_19_trfwwbasiccell_temp2_0: LUT4 
  generic map(
    INIT => X"C693"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(94),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(95),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_19_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_17x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(32),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(40),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_16x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(33),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(41),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_29x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(20),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(28),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_50_trfwwbasiccell_temp2_0: LUT4 
  generic map(
    INIT => X"C693"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(63),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_48_trfwwbasiccell_temp2_0: LUT4_L 
  generic map(
    INIT => X"C693"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(65),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_TEMP2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_49_trfwwbasiccell_temp2_1_0: LUT4_L 
  generic map(
    INIT => X"C693"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(65),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_TEMP2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_46x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(11),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_45x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(12),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_38x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(11),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_37x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(20),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_36x: LUT3 
  generic map(
    INIT => X"27"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(13),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_s_8_0_53x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TOPBITSIN(6),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(53));
  x_grlfpc2_0_r_i_pcce_2x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_V_I_EXEC_0_SQMUXA,
    I1 => holdn,
    O => N_5258);
  x_grlfpc2_0_comb_fpdecode_mov5: LUT3 
  generic map(
    INIT => X"40"
  )
  port map (
    I0 => cpi_d_inst(12),
    I1 => GRLFPC2_0_COMB_FPDECODE_MOV5_1,
    I2 => GRLFPC2_0_MOV_2_SQMUXA_1_0,
    O => GRLFPC2_0_COMB_FPDECODE_MOV5);
  x_grlfpc2_0_comb_un2_holdn: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_N_691,
    I1 => holdn,
    O => GRLFPC2_0_COMB_UN2_HOLDN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_12: LUT4 
  generic map(
    INIT => X"936C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1000,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_1(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_12_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_11: LUT4 
  generic map(
    INIT => X"936C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_999,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_1(11),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_11_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_10: LUT4 
  generic map(
    INIT => X"936C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_998,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_1(10),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_10_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_entryshft_un14_s_mov: LUT4 
  generic map(
    INIT => X"2A00"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN14_S_MOV_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(79),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(83),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN14_S_MOV);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_wqstsets_1_5x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN5_NOTAZERODENORM_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_4(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_5(5),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2002);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_aebeexc_un37_notbinfnan: LUT4_L 
  generic map(
    INIT => X"C080"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN11_NOTBINFNAN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTBINFNAN_4,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTBINFNAN_5,
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP1,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTBINFNAN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_aebeexc_un37_notainfnan: LUT4_L 
  generic map(
    INIT => X"C080"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN11_NOTAINFNAN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTAINFNAN_4,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTAINFNAN_5,
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP1,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTAINFNAN);
  x_grlfpc2_0_mov_7_sqmuxa: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => cpi_d_inst(19),
    I1 => GRLFPC2_0_COMB_FPDECODE_AFQ12,
    I2 => GRLFPC2_0_COMB_FPDECODE_UN3_OP,
    O => GRLFPC2_0_MOV_7_SQMUXA);
  x_grlfpc2_0_comb_fpdecode_rs2d5: LUT3 
  generic map(
    INIT => X"40"
  )
  port map (
    I0 => cpi_d_inst(12),
    I1 => GRLFPC2_0_COMB_FPDECODE_RS2D5_1,
    I2 => GRLFPC2_0_COMB_FPDECODE_RS2D5_3,
    O => GRLFPC2_0_COMB_FPDECODE_RS2D5);
  x_grlfpc2_0_comb_un6_iuexec: LUT4 
  generic map(
    INIT => X"0400"
  )
  port map (
    I0 => GRLFPC2_0_N_777,
    I1 => GRLFPC2_0_N_782,
    I2 => GRLFPC2_0_R_MK_BUSY,
    I3 => GRLFPC2_0_R_MK_BUSY2,
    O => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_wren2_2_sqmuxa: LUT4 
  generic map(
    INIT => X"1000"
  )
  port map (
    I0 => cpi_x_inst(20),
    I1 => GRLFPC2_0_R_X_AFSR,
    I2 => GRLFPC2_0_R_X_LD,
    I3 => GRLFPC2_0_WREN2_1_SQMUXA_1,
    O => GRLFPC2_0_WREN2_2_SQMUXA);
  x_grlfpc2_0_comb_fpdecode_mov6: LUT4 
  generic map(
    INIT => X"2000"
  )
  port map (
    I0 => cpi_d_inst(5),
    I1 => cpi_d_inst(6),
    I2 => GRLFPC2_0_COMB_FPDECODE_MOV6_2,
    I3 => GRLFPC2_0_MOV_2_SQMUXA_1_1,
    O => GRLFPC2_0_COMB_FPDECODE_MOV6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlaregxz_un7_xzaregloaden: LUT4 
  generic map(
    INIT => X"0002"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(6),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2023);
  x_grlfpc2_0_mov_5_sqmuxa_2: LUT4 
  generic map(
    INIT => X"4000"
  )
  port map (
    I0 => cpi_d_inst(10),
    I1 => GRLFPC2_0_COMB_FPDECODE_AFQ12,
    I2 => GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_1_0,
    I3 => GRLFPC2_0_MOV_2_SQMUXA_2,
    O => GRLFPC2_0_MOV_5_SQMUXA_2);
  x_grlfpc2_0_mov_0_sqmuxa_2_0: LUT4 
  generic map(
    INIT => X"2000"
  )
  port map (
    I0 => cpi_d_inst(12),
    I1 => cpi_d_inst(30),
    I2 => GRLFPC2_0_COMB_FPDECODE_MOV5_1,
    I3 => GRLFPC2_0_MOV_0_SQMUXA_3,
    O => GRLFPC2_0_MOV_0_SQMUXA_2_0);
  x_grlfpc2_0_v_state_1_sqmuxa_3_0: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_R_X_AFQ,
    I1 => GRLFPC2_0_SEQERR_1_SQMUXA_1_SN,
    I2 => GRLFPC2_0_WREN2_1_SQMUXA_1,
    O => GRLFPC2_0_V_STATE_1_SQMUXA_3_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_entryshft_entrypoint_0: LUT4_L 
  generic map(
    INIT => X"1555"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_S_CMP,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_ENTRYSHFT_S_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(82),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_0,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_ENTRYPOINT_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_waitmulxff_notsampledwait_0: LUT4 
  generic map(
    INIT => X"8A88"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CONDMUXMULXFF_UN4_NOTSQRTLFTCC,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(44),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_14_m_0_171x: LUT4 
  generic map(
    INIT => X"EE15"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(374),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(375),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(376),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(377),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14_M_0(171));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un79_zero: LUT3 
  generic map(
    INIT => X"7E"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(8),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un9_notprop: LUT2_L 
  generic map(
    INIT => X"6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(2),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN9_NOTPROP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un31_zero: LUT3 
  generic map(
    INIT => X"7E"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un55_zero: LUT3 
  generic map(
    INIT => X"7E"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(4),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_multiplelogic_un8_zero: LUT3 
  generic map(
    INIT => X"7E"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO);
  x_grlfpc2_0_comb_v_fsr_nonstd_1_m1_0_0: LUT3_L 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(22),
    I1 => GRLFPC2_0_R_FSR_NONSTD,
    I2 => GRLFPC2_0_V_FSR_AEXC_1_SQMUXA_SN,
    LO => GRLFPC2_0_COMB_V_FSR_NONSTD_1_M1);
  x_grlfpc2_0_comb_v_fsr_rd_1_m1_0_1x: LUT3_L 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(31),
    I1 => GRLFPC2_0_R_FSR_RD(1),
    I2 => GRLFPC2_0_V_FSR_AEXC_1_SQMUXA_SN,
    LO => GRLFPC2_0_COMB_V_FSR_RD_1_M1(1));
  x_grlfpc2_0_comb_v_fsr_rd_1_m1_0_0x: LUT3_L 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(30),
    I1 => GRLFPC2_0_R_FSR_RD(0),
    I2 => GRLFPC2_0_V_FSR_AEXC_1_SQMUXA_SN,
    LO => GRLFPC2_0_COMB_V_FSR_RD_1_M1(0));
  x_grlfpc2_0_comb_v_fsr_tem_1_m1_0_4x: LUT3_L 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(27),
    I1 => GRLFPC2_0_R_FSR_TEM(4),
    I2 => GRLFPC2_0_V_FSR_AEXC_1_SQMUXA_SN,
    LO => GRLFPC2_0_COMB_V_FSR_TEM_1_M1(4));
  x_grlfpc2_0_comb_v_fsr_tem_1_m1_0_3x: LUT3_L 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(26),
    I1 => GRLFPC2_0_R_FSR_TEM(3),
    I2 => GRLFPC2_0_V_FSR_AEXC_1_SQMUXA_SN,
    LO => GRLFPC2_0_COMB_V_FSR_TEM_1_M1(3));
  x_grlfpc2_0_comb_v_fsr_tem_1_m1_0_2x: LUT3_L 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(25),
    I1 => GRLFPC2_0_R_FSR_TEM(2),
    I2 => GRLFPC2_0_V_FSR_AEXC_1_SQMUXA_SN,
    LO => GRLFPC2_0_COMB_V_FSR_TEM_1_M1(2));
  x_grlfpc2_0_comb_v_fsr_tem_1_m1_0_1x: LUT3_L 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(24),
    I1 => GRLFPC2_0_R_FSR_TEM(1),
    I2 => GRLFPC2_0_V_FSR_AEXC_1_SQMUXA_SN,
    LO => GRLFPC2_0_COMB_V_FSR_TEM_1_M1(1));
  x_grlfpc2_0_comb_v_fsr_tem_1_m1_0_0x: LUT3_L 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(23),
    I1 => GRLFPC2_0_R_FSR_TEM(0),
    I2 => GRLFPC2_0_V_FSR_AEXC_1_SQMUXA_SN,
    LO => GRLFPC2_0_COMB_V_FSR_TEM_1_M1(0));
  x_grlfpc2_0_comb_v_fsr_fcc_1_m0_0_1x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(11),
    I1 => CPO_CC_1_INT_4,
    I2 => GRLFPC2_0_V_FSR_AEXC_1_SQMUXA_SN,
    O => GRLFPC2_0_COMB_V_FSR_FCC_1_M0(1));
  x_grlfpc2_0_comb_v_fsr_fcc_1_m0_0_0x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(10),
    I1 => CPO_CC_0_INT_3,
    I2 => GRLFPC2_0_V_FSR_AEXC_1_SQMUXA_SN,
    O => GRLFPC2_0_COMB_V_FSR_FCC_1_M0(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_ss12_0: LUT4 
  generic map(
    INIT => X"7F55"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_53_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SM3_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV_4_0,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV_6_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SS12);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un4_temp_u_0_0x: LUT4 
  generic map(
    INIT => X"80BF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_104,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_16_REP1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(5),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN4_TEMP(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_7x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(49),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(224),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_114);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_8x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(48),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(223),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_115);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_9x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(47),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(222),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_116);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_10x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(46),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(221),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_117);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_11x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(45),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(220),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_118);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_12x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(44),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(219),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_119);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_13x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(43),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(218),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_120);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_14x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(217),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_121);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_15x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(41),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(216),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_122);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_16x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(215),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_123);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_18x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(38),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(213),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_125);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_19x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(37),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(212),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_126);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_20x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(36),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(211),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_127);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_21x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(35),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(210),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_128);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_22x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(34),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(209),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_129);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_25x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(31),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(206),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_132);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_26x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(205),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_133);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_27x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(204),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_134);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_28x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(28),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(203),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_135);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_30x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(26),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(201),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_137);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_31x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(25),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(200),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_138);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_32x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(24),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(199),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_139);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_33x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(198),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_140);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_34x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(22),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(197),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_141);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_35x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(196),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_142);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_36x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(20),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(195),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_143);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_37x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(194),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_144);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_38x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(18),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(193),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_145);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_39x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(192),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_146);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_40x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(191),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_147);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_41x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(15),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(190),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_148);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_42x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(14),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(189),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_149);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_43x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(13),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(188),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_150);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_47x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(9),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(184),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_154);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_49x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(182),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_156);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_50x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(181),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_157);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_51x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(180),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_158);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_52x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(179),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_159);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_54x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(177),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_161);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_55x: LUT4 
  generic map(
    INIT => X"ECE4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(176),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(10),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_162);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_am_0x: LUT4 
  generic map(
    INIT => X"B0F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP1,
    O => N_12094);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_bm_0x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(244),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(257),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
    O => N_12095);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_0x: MUXF5 port map (
      I0 => N_12094,
      I1 => N_12095,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_am_1x: LUT4 
  generic map(
    INIT => X"E0A0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP1,
    O => N_12096);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_bm_1x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(243),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(256),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
    O => N_12097);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_1x: MUXF5 port map (
      I0 => N_12096,
      I1 => N_12097,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_am_3x: LUT4 
  generic map(
    INIT => X"A0E0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP1,
    O => N_12098);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_bm_3x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(241),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(254),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
    O => N_12099);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_3x: MUXF5 port map (
      I0 => N_12098,
      I1 => N_12099,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_am_7x: LUT4 
  generic map(
    INIT => X"0080"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP1,
    O => N_12100);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_bm_7x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(237),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(250),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
    O => N_12101);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_7x: MUXF5 port map (
      I0 => N_12100,
      I1 => N_12101,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_am_8x: LUT4 
  generic map(
    INIT => X"0080"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP1,
    O => N_12102);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_bm_8x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(236),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(249),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
    O => N_12103);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_8x: MUXF5 port map (
      I0 => N_12102,
      I1 => N_12103,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_am_9x: LUT4 
  generic map(
    INIT => X"0080"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP1,
    O => N_12104);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_bm_9x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(235),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(248),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
    O => N_12105);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_expxbus_3_0_9x: MUXF5 port map (
      I0 => N_12104,
      I1 => N_12105,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(9));
  x_grlfpc2_0_op1_0_32x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(0),
    I2 => rfo2_data1(0),
    O => GRLFPC2_0_OP1(32));
  x_grlfpc2_0_op1_0_33x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(1),
    I2 => rfo2_data1(1),
    O => GRLFPC2_0_OP1(33));
  x_grlfpc2_0_op1_0_34x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(2),
    I2 => rfo2_data1(2),
    O => GRLFPC2_0_OP1(34));
  x_grlfpc2_0_op1_0_35x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(3),
    I2 => rfo2_data1(3),
    O => GRLFPC2_0_OP1(35));
  x_grlfpc2_0_op1_0_36x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(4),
    I2 => rfo2_data1(4),
    O => GRLFPC2_0_OP1(36));
  x_grlfpc2_0_op1_0_37x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(5),
    I2 => rfo2_data1(5),
    O => GRLFPC2_0_OP1(37));
  x_grlfpc2_0_op1_0_38x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(6),
    I2 => rfo2_data1(6),
    O => GRLFPC2_0_OP1(38));
  x_grlfpc2_0_op1_0_39x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(7),
    I2 => rfo2_data1(7),
    O => GRLFPC2_0_OP1(39));
  x_grlfpc2_0_op1_0_40x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(8),
    I2 => rfo2_data1(8),
    O => GRLFPC2_0_OP1(40));
  x_grlfpc2_0_op1_0_41x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(9),
    I2 => rfo2_data1(9),
    O => GRLFPC2_0_OP1(41));
  x_grlfpc2_0_op1_0_42x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(10),
    I2 => rfo2_data1(10),
    O => GRLFPC2_0_OP1(42));
  x_grlfpc2_0_op1_0_43x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(11),
    I2 => rfo2_data1(11),
    O => GRLFPC2_0_OP1(43));
  x_grlfpc2_0_op1_0_47x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(15),
    I2 => rfo2_data1(15),
    O => GRLFPC2_0_OP1(47));
  x_grlfpc2_0_op1_0_49x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(17),
    I2 => rfo2_data1(17),
    O => GRLFPC2_0_OP1(49));
  x_grlfpc2_0_op1_0_51x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(19),
    I2 => rfo2_data1(19),
    O => GRLFPC2_0_OP1(51));
  x_grlfpc2_0_op1_0_52x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(20),
    I2 => rfo2_data1(20),
    O => GRLFPC2_0_OP1(52));
  x_grlfpc2_0_op1_0_55x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(23),
    I2 => rfo2_data1(23),
    O => GRLFPC2_0_OP1(55));
  x_grlfpc2_0_op1_0_56x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(24),
    I2 => rfo2_data1(24),
    O => GRLFPC2_0_OP1(56));
  x_grlfpc2_0_op1_0_59x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(27),
    I2 => rfo2_data1(27),
    O => GRLFPC2_0_OP1(59));
  x_grlfpc2_0_op1_0_62x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(30),
    I2 => rfo2_data1(30),
    O => GRLFPC2_0_OP1(62));
  x_grlfpc2_0_op1_0_63x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(31),
    I2 => rfo2_data1(31),
    O => GRLFPC2_0_OP1(63));
  x_grlfpc2_0_op2_0_32x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(0),
    I2 => rfo2_data2(0),
    O => GRLFPC2_0_OP2(32));
  x_grlfpc2_0_op2_0_33x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(1),
    I2 => rfo2_data2(1),
    O => GRLFPC2_0_OP2(33));
  x_grlfpc2_0_op2_0_34x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(2),
    I2 => rfo2_data2(2),
    O => GRLFPC2_0_OP2(34));
  x_grlfpc2_0_op2_0_35x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(3),
    I2 => rfo2_data2(3),
    O => GRLFPC2_0_OP2(35));
  x_grlfpc2_0_op2_0_36x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(4),
    I2 => rfo2_data2(4),
    O => GRLFPC2_0_OP2(36));
  x_grlfpc2_0_op2_0_37x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(5),
    I2 => rfo2_data2(5),
    O => GRLFPC2_0_OP2(37));
  x_grlfpc2_0_op2_0_38x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(6),
    I2 => rfo2_data2(6),
    O => GRLFPC2_0_OP2(38));
  x_grlfpc2_0_op2_0_39x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(7),
    I2 => rfo2_data2(7),
    O => GRLFPC2_0_OP2(39));
  x_grlfpc2_0_op2_0_40x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(8),
    I2 => rfo2_data2(8),
    O => GRLFPC2_0_OP2(40));
  x_grlfpc2_0_op2_0_41x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(9),
    I2 => rfo2_data2(9),
    O => GRLFPC2_0_OP2(41));
  x_grlfpc2_0_op2_0_42x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(10),
    I2 => rfo2_data2(10),
    O => GRLFPC2_0_OP2(42));
  x_grlfpc2_0_op2_0_44x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(12),
    I2 => rfo2_data2(12),
    O => GRLFPC2_0_OP2(44));
  x_grlfpc2_0_op2_0_45x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(13),
    I2 => rfo2_data2(13),
    O => GRLFPC2_0_OP2(45));
  x_grlfpc2_0_op2_0_47x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(15),
    I2 => rfo2_data2(15),
    O => GRLFPC2_0_OP2(47));
  x_grlfpc2_0_op2_0_48x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(16),
    I2 => rfo2_data2(16),
    O => GRLFPC2_0_OP2(48));
  x_grlfpc2_0_op2_0_49x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(17),
    I2 => rfo2_data2(17),
    O => GRLFPC2_0_OP2(49));
  x_grlfpc2_0_op2_0_50x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(18),
    I2 => rfo2_data2(18),
    O => GRLFPC2_0_OP2(50));
  x_grlfpc2_0_op2_0_51x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(19),
    I2 => rfo2_data2(19),
    O => GRLFPC2_0_OP2(51));
  x_grlfpc2_0_op2_0_52x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(20),
    I2 => rfo2_data2(20),
    O => GRLFPC2_0_OP2(52));
  x_grlfpc2_0_op2_0_53x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(21),
    I2 => rfo2_data2(21),
    O => GRLFPC2_0_OP2(53));
  x_grlfpc2_0_op2_0_55x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(23),
    I2 => rfo2_data2(23),
    O => GRLFPC2_0_OP2(55));
  x_grlfpc2_0_op2_0_56x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(24),
    I2 => rfo2_data2(24),
    O => GRLFPC2_0_OP2(56));
  x_grlfpc2_0_op2_0_57x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(25),
    I2 => rfo2_data2(25),
    O => GRLFPC2_0_OP2(57));
  x_grlfpc2_0_op2_0_58x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(26),
    I2 => rfo2_data2(26),
    O => GRLFPC2_0_OP2(58));
  x_grlfpc2_0_op2_0_59x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(27),
    I2 => rfo2_data2(27),
    O => GRLFPC2_0_OP2(59));
  x_grlfpc2_0_op2_0_60x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(28),
    I2 => rfo2_data2(28),
    O => GRLFPC2_0_OP2(60));
  x_grlfpc2_0_op2_0_61x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(29),
    I2 => rfo2_data2(29),
    O => GRLFPC2_0_OP2(61));
  x_grlfpc2_0_op2_0_62x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(30),
    I2 => rfo2_data2(30),
    O => GRLFPC2_0_OP2(62));
  x_grlfpc2_0_op2_0_63x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(31),
    I2 => rfo2_data2(31),
    O => GRLFPC2_0_OP2(63));
  x_grlfpc2_0_wrdata_0_0_63x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(31),
    I1 => GRLFPC2_0_R_I_RES(63),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_126);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_48x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(183),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_155);
  x_grlfpc2_0_op1_0_46x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(14),
    I2 => rfo2_data1(14),
    O => GRLFPC2_0_OP1(46));
  x_grlfpc2_0_op1_0_45x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(13),
    I2 => rfo2_data1(13),
    O => GRLFPC2_0_OP1(45));
  x_grlfpc2_0_op1_0_58x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(26),
    I2 => rfo2_data1(26),
    O => GRLFPC2_0_OP1(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m12_0_am_0x: LUT3 
  generic map(
    INIT => X"BA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5),
    O => N_12106);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m12_0_bm_0x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SM3_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(11),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(13),
    LO => N_12107);
  x_grlfpc2_0_op1_0_61x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(29),
    I2 => rfo2_data1(29),
    O => GRLFPC2_0_OP1(61));
  x_grlfpc2_0_op1_0_60x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(28),
    I2 => rfo2_data1(28),
    O => GRLFPC2_0_OP1(60));
  x_grlfpc2_0_op1_0_57x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(25),
    I2 => rfo2_data1(25),
    O => GRLFPC2_0_OP1(57));
  x_grlfpc2_0_I_189_0_am: LUT2 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => cpi_d_inst(25),
    I1 => GRLFPC2_0_MOV_7_SQMUXA_3,
    O => N_12108);
  x_grlfpc2_0_I_189_0_bm: LUT3 
  generic map(
    INIT => X"20"
  )
  port map (
    I0 => cpi_d_inst(20),
    I1 => cpi_d_inst(22),
    I2 => GRLFPC2_0_N_703_1,
    O => N_12109);
  x_grlfpc2_0_I_189_0: MUXF5 port map (
      I0 => N_12108,
      I1 => N_12109,
      S => cpi_d_inst(19),
      O => GRLFPC2_0_N_634);
  x_grlfpc2_0_op1_0_48x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(16),
    I2 => rfo2_data1(16),
    O => GRLFPC2_0_OP1(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_56x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(175),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_163);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_46x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(10),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(185),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_153);
  x_grlfpc2_0_op2_0_43x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(11),
    I2 => rfo2_data2(11),
    O => GRLFPC2_0_OP2(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_6x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(50),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(225),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_113);
  x_grlfpc2_0_op2_0_46x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(14),
    I2 => rfo2_data2(14),
    O => GRLFPC2_0_OP2(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_17x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(214),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_124);
  x_grlfpc2_0_op2_0_54x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(22),
    I2 => rfo2_data2(22),
    O => GRLFPC2_0_OP2(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_24x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(32),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(207),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_131);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_23x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(33),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(208),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_130);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_29x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(27),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(202),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_136);
  x_grlfpc2_0_op1_0_54x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(22),
    I2 => rfo2_data1(22),
    O => GRLFPC2_0_OP1(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_44x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(187),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_151);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_53x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(178),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_160);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_45x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(11),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(186),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_152);
  x_grlfpc2_0_op1_0_53x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(21),
    I2 => rfo2_data1(21),
    O => GRLFPC2_0_OP1(53));
  x_grlfpc2_0_op1_0_50x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(18),
    I2 => rfo2_data1(18),
    O => GRLFPC2_0_OP1(50));
  x_grlfpc2_0_op1_0_44x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_772,
    I1 => rfo1_data1(12),
    I2 => rfo2_data1(12),
    O => GRLFPC2_0_OP1(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_si_114_1_1_0_56x: LUT3 
  generic map(
    INIT => X"A6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(57),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(316),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_114_1_1_0(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_5_sqmuxa_2: LUT3 
  generic map(
    INIT => X"20"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_3_sqmuxa_2_1: LUT3 
  generic map(
    INIT => X"08"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_un57_shdvar: LUT4 
  generic map(
    INIT => X"7F00"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_NOTAM2_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_6_AND_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_7_AND1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(3),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN57_SHDVAR);
  x_grlfpc2_0_un1_fpci_5: LUT4 
  generic map(
    INIT => X"08AA"
  )
  port map (
    I0 => GRLFPC2_0_N_781,
    I1 => GRLFPC2_0_R_X_AFSR,
    I2 => GRLFPC2_0_R_X_LD,
    I3 => GRLFPC2_0_V_STATE_1_SQMUXA_1,
    O => GRLFPC2_0_N_755);
  x_grlfpc2_0_I_204: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_FPDECODE_RS2D5,
    I1 => GRLFPC2_0_MOV_7_SQMUXA,
    O => GRLFPC2_0_N_653);
  x_grlfpc2_0_comb_v_a_afsr_1s2_279: LUT4 
  generic map(
    INIT => X"0E0F"
  )
  port map (
    I0 => cpi_d_inst(19),
    I1 => cpi_d_inst(23),
    I2 => GRLFPC2_0_COMB_FPDECODE_AFQ3,
    I3 => GRLFPC2_0_MOV_7_SQMUXA_3,
    O => GRLFPC2_0_RS1V10_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus24: LUT3 
  generic map(
    INIT => X"20"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTXZYFROMD_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24);
  x_grlfpc2_0_comb_rs2_1_sn_m1: LUT2 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => GRLFPC2_0_RS2_0_SQMUXA,
    I1 => holdn,
    O => GRLFPC2_0_COMB_RS2_1_SN_N_2);
  x_grlfpc2_0_comb_seqerr_un13_op: LUT4 
  generic map(
    INIT => X"DC00"
  )
  port map (
    I0 => cpi_d_inst(23),
    I1 => GRLFPC2_0_COMB_FPDECODE_AFQ7,
    I2 => GRLFPC2_0_COMB_FPDECODE_AFQ8_0,
    I3 => GRLFPC2_0_COMB_FPDECODE_AFQ13,
    O => GRLFPC2_0_COMB_SEQERR_UN13_OP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_Excep_1_0x: LUT4 
  generic map(
    INIT => X"FAEE"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2003,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN3_INEXACT,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT,
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1990);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m13_0_am_1x: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SM6_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SS6,
    O => N_12110);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m13_0_bm_1x: LUT3 
  generic map(
    INIT => X"B1"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SM0_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(15),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
    O => N_12111);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m13_0_1x: MUXF5 port map (
      I0 => N_12110,
      I1 => N_12111,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV_6,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M13(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m13_0_am_2x: LUT2 
  generic map(
    INIT => X"D"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SM6_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SS6,
    O => N_12112);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m13_0_bm_2x: LUT2 
  generic map(
    INIT => X"D"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SM0_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
    O => N_12113);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m13_0_2x: MUXF5 port map (
      I0 => N_12112,
      I1 => N_12113,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV_6,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M13(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m12_0_am_1x: LUT3 
  generic map(
    INIT => X"54"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5),
    O => N_12114);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m12_0_bm_1x: LUT3 
  generic map(
    INIT => X"B1"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SM3_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(11),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(13),
    O => N_12115);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m12_0_1x: MUXF5 port map (
      I0 => N_12114,
      I1 => N_12115,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV_6,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M12(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m12_0_am_2x: LUT3 
  generic map(
    INIT => X"01"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5),
    O => N_12116);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m12_0_bm_2x: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SM3_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(13),
    O => N_12117);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m12_0_2x: MUXF5 port map (
      I0 => N_12116,
      I1 => N_12117,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV_6,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M12(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_7_0_0_am: LUT3 
  generic map(
    INIT => X"95"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(48),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(52),
    I2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => N_12118);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_7_0_0_bm: LUT4 
  generic map(
    INIT => X"A5C3"
  )
  port map (
    I0 => N_2477,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_AREGXORBREG,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(48),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(52),
    O => N_12119);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_7_0_0: MUXF5 port map (
      I0 => N_12118,
      I1 => N_12119,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(51),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_353);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m13_0_0x: LUT4 
  generic map(
    INIT => X"D8F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_53_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M2(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SS6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV_6_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M13(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_wqsctrl_1_68x: LUT4 
  generic map(
    INIT => X"4000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(12),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_2_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(47),
    I3 => rst,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_1(68));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_wqstsets_1_4x: LUT4 
  generic map(
    INIT => X"0203"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN5_NOTBZERODENORM_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTBINFNAN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(246),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_wqstsets_1_3x: LUT4 
  generic map(
    INIT => X"0203"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN5_NOTAZERODENORM_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN37_NOTAINFNAN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(233),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un17_wqstsets: LUT4 
  generic map(
    INIT => X"1101"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1991,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN5_NOTSHIFTCOUNT1_0,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN17_WQSTSETS);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_temp_1: LUT4 
  generic map(
    INIT => X"0100"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN14_S_MOV,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN23_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(73),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP_1);
  x_grlfpc2_0_afq_3_sqmuxa: LUT4 
  generic map(
    INIT => X"4000"
  )
  port map (
    I0 => cpi_d_inst(19),
    I1 => cpi_d_inst(20),
    I2 => GRLFPC2_0_COMB_FPDECODE_AFQ4_1,
    I3 => GRLFPC2_0_COMB_FPDECODE_AFQ13,
    O => GRLFPC2_0_AFQ_3_SQMUXA);
  x_grlfpc2_0_comb_un8_ccv: LUT4 
  generic map(
    INIT => X"0222"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN8_CCV_1,
    I1 => GRLFPC2_0_COMB_UN14_CCV,
    I2 => GRLFPC2_0_R_I_EXEC,
    I3 => GRLFPC2_0_R_I_INST(19),
    O => cpo_ccv);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus25: LUT3 
  generic map(
    INIT => X"40"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTXZYFROMD_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus26: LUT3 
  generic map(
    INIT => X"08"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTXZYFROMD_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26);
  x_grlfpc2_0_wren2_1_sqmuxa_1_0: LUT4 
  generic map(
    INIT => X"2000"
  )
  port map (
    I0 => cpi_x_inst(20),
    I1 => GRLFPC2_0_R_X_AFSR,
    I2 => GRLFPC2_0_R_X_LD,
    I3 => GRLFPC2_0_WREN2_1_SQMUXA_1,
    O => GRLFPC2_0_WREN2_1_SQMUXA_1_0);
  x_grlfpc2_0_comb_fpdecode_un1_wren210: LUT4 
  generic map(
    INIT => X"4000"
  )
  port map (
    I0 => cpi_d_inst(7),
    I1 => cpi_d_inst(12),
    I2 => GRLFPC2_0_COMB_FPDECODE_RS2D5_1,
    I3 => GRLFPC2_0_COMB_FPDECODE_RS2D5_3,
    O => GRLFPC2_0_COMB_FPDECODE_UN1_WREN210);
  x_grlfpc2_0_I_162_266_138_tz: LUT4_L 
  generic map(
    INIT => X"3011"
  )
  port map (
    I0 => GRLFPC2_0_ANNULFPU_0_SQMUXA_1,
    I1 => GRLFPC2_0_ANNULRES_0_SQMUXA_3_0,
    I2 => GRLFPC2_0_COMB_UN1_FPCI_1_I,
    I3 => GRLFPC2_0_R_M_FPOP,
    LO => N_2291_TZ);
  x_grlfpc2_0_comb_rsdecode_rs1v2_0: LUT4 
  generic map(
    INIT => X"2333"
  )
  port map (
    I0 => cpi_d_inst(12),
    I1 => GRLFPC2_0_COMB_FPDECODE_MOV6,
    I2 => GRLFPC2_0_COMB_FPDECODE_UN1_FPCI_1_0,
    I3 => GRLFPC2_0_MOV_0_SQMUXA_2,
    O => GRLFPC2_0_COMB_RSDECODE_RS1V2_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_2_1_0x: LUT4 
  generic map(
    INIT => X"0E00"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2030,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN46_XZYBUSLSBS,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_I(15),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_2_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_9_sqmuxa_m1_e_0: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA_M1_E_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_UN99_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_UN96_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_49_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"7E00"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(4),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_TEMP2_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_50_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_UN531_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_UN528_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_50_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_UN360_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_UN357_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_51_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_UN357_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_UN354_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_48_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"7E00"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(4),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_TEMP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_46_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_UN543_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_UN540_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_45_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_UN546_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_UN543_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_47_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_UN540_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_UN537_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_38_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_UN396_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_UN393_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_36_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_UN573_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_UN570_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_32_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_UN243_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_UN240_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_35_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_UN576_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_UN573_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_36_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_UN402_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_UN399_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_UN612_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_UN609_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_27_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_UN429_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_UN426_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_I_193: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => cpi_d_inst(30),
    I1 => GRLFPC2_0_N_634,
    O => GRLFPC2_0_N_635);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_13_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_UN129_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_UN126_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_UN660_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_UN657_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_12_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_UN132_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_UN129_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_13_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_UN300_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_UN297_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_13_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_UN471_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_UN468_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_14_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_UN468_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_UN465_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_UN135_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_UN132_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_27_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_UN87_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_UN84_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_1_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_UN678_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_UN675_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_UN675_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_UN672_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_UN672_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_UN669_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_UN159_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_UN156_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_1_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_UN165_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_UN162_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_0_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_UN168_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_UN165_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_1_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_UN336_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_UN333_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_34_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_UN237_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_UN234_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_15_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_UN123_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_UN120_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_16_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_UN291_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_UN288_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_15_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_UN294_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_UN291_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_14_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_UN297_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_UN294_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_UN312_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_UN309_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_25_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_UN264_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_UN261_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_21_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_UN105_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_UN102_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_16_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_UN462_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_UN459_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_19_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_19_TRFWWBASICCELL_UN111_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_UN108_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_19_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_15_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"7E00"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(4),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_TEMP2_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_21_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_UN447_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_UN444_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_49_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"7E00"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(2),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_TEMP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_49_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_UN534_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_UN531_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_UN441_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_UN438_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_22_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_UN444_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_UN441_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_20_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_UN450_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_UN447_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_48_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_UN366_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_UN363_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_49_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_UN363_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_UN360_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_47_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_UN369_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_UN366_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_14_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_UN126_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_UN123_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_8_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_UN315_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_UN312_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_UN348_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_UN345_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"160E"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(4),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(58),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_29_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_UN594_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_UN591_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_53_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_UN351_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_UN348_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_52_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_UN525_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_UN522_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_51_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_UN528_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_UN525_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_12_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_UN645_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_UN642_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_52_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_UN354_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_UN351_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_13_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_UN642_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_UN639_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_UN483_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_UN480_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_8_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_UN486_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_UN483_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_43_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_UN552_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_UN549_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_42_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_UN555_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_UN552_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_27_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_UN600_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_UN597_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_26_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_UN603_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_UN600_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_28_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_UN255_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_UN252_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_29_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_UN423_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_UN420_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_28_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_UN426_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_UN423_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_26_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_UN90_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_UN87_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_21_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_UN618_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_UN615_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_UN489_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_UN486_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_UN480_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_UN477_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_35_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_UN405_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_UN402_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_12_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_UN474_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_UN471_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_44_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_UN378_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_UN375_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_UN501_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_UN498_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_UN504_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_UN501_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_1_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_UN507_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_UN504_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_0_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_UN510_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_UN507_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_45_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_UN375_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_UN372_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_46_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_UN372_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_UN369_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_50_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_UN18_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_UN15_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_51_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_UN186_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_UN183_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_UN477_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_UN474_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_30_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_UN420_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_UN417_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_35_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_UN63_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_UN60_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_28_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_UN597_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_UN594_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_33_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_UN411_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_UN408_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_32_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_UN414_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_UN411_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_36_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_UN60_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_UN57_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_37_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_UN57_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_UN54_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_37_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_UN228_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_UN225_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_35_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_UN234_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_UN231_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_18_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_18_TRFWWBASICCELL_UN114_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_19_TRFWWBASICCELL_UN111_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_18_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_0_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_UN339_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_UN336_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_6_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_UN150_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_UN147_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_UN141_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_UN138_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_8_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_UN144_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_UN141_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_5_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_UN495_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_UN492_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_21_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_UN276_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_UN273_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_17_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_UN630_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_18_TRFWWBASICCELL_UN627_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_16_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_UN633_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_UN630_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_29_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_UN81_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_UN78_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_27_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_UN258_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_UN255_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_12_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_UN303_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_UN300_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_UN306_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_UN303_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"160E"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(4),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(58),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_55_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_UN174_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_UN171_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_UN6_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_UN3_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_53_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_UN9_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_UN6_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_5: LUT4_L 
  generic map(
    INIT => X"6C93"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1017,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_32_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_UN72_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_UN69_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_34_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_UN66_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_UN63_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_17_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_UN117_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_18_TRFWWBASICCELL_UN114_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_46_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"7E00"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(2),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_TEMP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_45_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_UN204_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_UN201_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_UN330_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_UN327_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_UN327_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_UN324_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_22_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_UN615_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_UN612_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_UN651_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_UN648_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_UN609_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_UN606_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_45_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_UN33_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_UN30_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_43_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_UN210_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_UN207_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"160E"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(2),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(58),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_UN438_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_UN435_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_46_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_UN201_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_UN198_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_25_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_UN93_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_UN90_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_22_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_UN102_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_UN99_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_55_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_UN3_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_28_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_UN84_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_UN81_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_UN654_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_UN651_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_UN648_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_UN645_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_39_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_UN51_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_UN48_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_39_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_UN222_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_UN219_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_UN318_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_UN315_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_48_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_UN537_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_UN534_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_53_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_UN522_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_UN519_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_UN519_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_UN516_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_55_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_UN516_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_UN513_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_UN138_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_UN135_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_6_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_UN492_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_UN489_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_19_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_19_TRFWWBASICCELL_UN624_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_UN621_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_19_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_52_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_UN12_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_UN9_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_33_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_UN240_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_UN237_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_47_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"7E00"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(2),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_TEMP2_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_41_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_UN558_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_UN555_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_15_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_UN636_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_UN633_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_6_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_UN321_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_UN318_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_41_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_UN45_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_UN42_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_32_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_UN585_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_UN582_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_44_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_UN207_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_UN204_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_25_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_UN435_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_UN432_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_26_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_UN432_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_UN429_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_UN309_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_UN306_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_31_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_UN417_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_UN414_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_34_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_UN408_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_UN405_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_37_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_UN399_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_UN396_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_39_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_UN393_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_UN390_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_40_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_UN390_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_UN387_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_41_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_UN387_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_UN384_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_42_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_UN384_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_UN381_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_43_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_UN381_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_UN378_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_48_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"7E00"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(2),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_TEMP2_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_UN498_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_UN495_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_20_trfwwbasiccell_cin_3: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_UN621_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_UN618_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_CIN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_34_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_UN579_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_UN576_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_51_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_UN15_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_UN12_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_20_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_UN108_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_UN105_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_30_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_UN78_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_UN75_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_22_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_UN273_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_UN270_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_UN270_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_UN267_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_UN267_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_UN264_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_26_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_UN261_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_UN258_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_44_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_UN549_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_UN546_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_33_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_UN582_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_UN579_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_UN96_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_UN93_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_25_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_UN606_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_UN603_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_30_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_UN591_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_UN588_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_43_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_UN39_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_UN36_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_33_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_UN69_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_UN66_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_52_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_UN183_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_UN180_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_53_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_UN180_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_UN177_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_UN177_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_UN174_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_UN162_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_UN159_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_UN156_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_UN153_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_5_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_UN153_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_UN150_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_UN147_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_UN144_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_36_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_UN231_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_UN228_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_40_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_UN48_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_UN45_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_38_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_UN225_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_UN222_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_42_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_UN42_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_UN39_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_UN333_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_UN330_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_31_trfwwbasiccell_cin_2: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_UN75_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_UN72_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_CIN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_5_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_UN324_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_UN321_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_18_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_18_TRFWWBASICCELL_UN627_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_19_TRFWWBASICCELL_UN624_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_18_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_40_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_UN219_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_UN216_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_31_trfwwbasiccell_cin_1: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_UN588_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_UN585_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_CIN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_38_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_UN54_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_UN51_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_8_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_UN657_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_UN654_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_6_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_UN663_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_UN660_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_44_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_UN36_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_UN33_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_55_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_3(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_UN345_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_UN342_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_40_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_UN561_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_UN558_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_UN669_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_UN666_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_14_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_UN639_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_UN636_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_31_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_2(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_UN246_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_UN243_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_5_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SHIFT(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_UN666_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_UN663_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_16_trfwwbasiccell_cin: LUT4 
  generic map(
    INIT => X"C840"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_SHIFT_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN8_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_UN120_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_UN117_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_CIN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_6x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(10),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_8x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_11x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(11),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(15),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_15x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(15),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(19),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_19x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(19),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(23),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_20x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(20),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(24),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_22x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(22),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(26),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_23x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(27),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_24x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(24),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(28),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_26x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(26),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_36x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(36),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_37x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(37),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(41),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_40x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(40),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(44),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_44x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(44),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(48),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_45x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(45),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(49),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_46x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(46),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(50),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_48x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(48),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(52),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_49x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(49),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_51x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(51),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_53x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(53),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(57),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_54x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(54),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(57),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_55x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(55),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(57),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_56x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(56),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(57),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(56));
  x_grlfpc2_0_comb_wraddr_5_0_2x: LUT4 
  generic map(
    INIT => X"AAB8"
  )
  port map (
    I0 => cpi_x_inst(27),
    I1 => GRLFPC2_0_COMB_UN1_R_I_V,
    I2 => GRLFPC2_0_R_I_INST(27),
    I3 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_COMB_WRADDR_5(2));
  x_grlfpc2_0_comb_wraddr_5_0_3x: LUT4 
  generic map(
    INIT => X"AAB8"
  )
  port map (
    I0 => cpi_x_inst(28),
    I1 => GRLFPC2_0_COMB_UN1_R_I_V,
    I2 => GRLFPC2_0_R_I_INST(28),
    I3 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_COMB_WRADDR_5(3));
  x_grlfpc2_0_comb_wraddr_5_0_4x: LUT4 
  generic map(
    INIT => X"AAB8"
  )
  port map (
    I0 => cpi_x_inst(29),
    I1 => GRLFPC2_0_COMB_UN1_R_I_V,
    I2 => GRLFPC2_0_R_I_INST(29),
    I3 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_COMB_WRADDR_5(4));
  x_grlfpc2_0_comb_rdd_3_0: LUT4 
  generic map(
    INIT => X"E4CC"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN1_R_I_V,
    I1 => GRLFPC2_0_R_I_RDD,
    I2 => GRLFPC2_0_R_X_RDD,
    I3 => GRLFPC2_0_V_I_EXEC_0_SQMUXA,
    O => GRLFPC2_0_COMB_RDD_3);
  x_grlfpc2_0_comb_wraddr_5_0_1x: LUT4 
  generic map(
    INIT => X"AAB8"
  )
  port map (
    I0 => cpi_x_inst(26),
    I1 => GRLFPC2_0_COMB_UN1_R_I_V,
    I2 => GRLFPC2_0_R_I_INST(26),
    I3 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_COMB_WRADDR_5(1));
  x_grlfpc2_0_comb_wraddr_5_0_0x: LUT4 
  generic map(
    INIT => X"AAB8"
  )
  port map (
    I0 => cpi_x_inst(25),
    I1 => GRLFPC2_0_COMB_UN1_R_I_V,
    I2 => GRLFPC2_0_R_I_INST(25),
    I3 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_COMB_WRADDR_5(0));
  x_grlfpc2_0_I_225_0: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => cpi_d_inst(19),
    I1 => GRLFPC2_0_COMB_FPDECODE_MOV5,
    I2 => GRLFPC2_0_COMB_FPDECODE_RS2D5,
    O => GRLFPC2_0_N_673);
  x_grlfpc2_0_comb_rs1d_1_m1_0_0: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => cpi_d_inst(20),
    I1 => GRLFPC2_0_COMB_FPDECODE_RS2D5,
    I2 => GRLFPC2_0_MOV_7_SQMUXA,
    O => GRLFPC2_0_COMB_RS1D_1_M1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_1x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_sn_m3_0: LUT3 
  generic map(
    INIT => X"68"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTXZYFROMD_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_21x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(25),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_17x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(17),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(21),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_13x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(13),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_47x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(47),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_43x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(43),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(47),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_42x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(42),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(46),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_39x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(39),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(43),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_38x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(38),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_4_2_0_41x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(41),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(45),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(41));
  x_grlfpc2_0_comb_annulfpu_1_u: LUT4 
  generic map(
    INIT => X"4044"
  )
  port map (
    I0 => GRLFPC2_0_N_206,
    I1 => GRLFPC2_0_COMB_ANNULFPU_1_U_0,
    I2 => GRLFPC2_0_COMB_UN1_FPCI_1_I,
    I3 => GRLFPC2_0_R_M_FPOP,
    O => GRLFPC2_0_N_710);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_NE_0: LUT4 
  generic map(
    INIT => X"8448"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(4),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_10_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_1(4),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_NE_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_1_41x: LUT4 
  generic map(
    INIT => X"2000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTXZYFROMD_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(41),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_1(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_1_39x: LUT4 
  generic map(
    INIT => X"2000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTXZYFROMD_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(39),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_1(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_3x: LUT4 
  generic map(
    INIT => X"2000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTXZYFROMD_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_174x: LUT4 
  generic map(
    INIT => X"0800"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTXZYFROMD_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(174),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(174));
  x_grlfpc2_0_mov_3_sqmuxa_1: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_COMB_FPDECODE_AFQ12,
    I1 => GRLFPC2_0_COMB_FPDECODE_MOV5,
    I2 => GRLFPC2_0_COMB_FPDECODE_MOV11,
    O => GRLFPC2_0_MOV_3_SQMUXA_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_oprexcshft_un3_oprexc: LUT4 
  generic map(
    INIT => X"4CCC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_AEBEEXC_UN5_NOTBZERODENORM_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_4(6),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_5(6),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_OPREXCSHFT_UN3_OPREXC);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un42_conditional: LUT2 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2002,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1(3),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN42_CONDITIONAL);
  x_grlfpc2_0_comb_fpdecode_mov3: LUT4 
  generic map(
    INIT => X"1333"
  )
  port map (
    I0 => GRLFPC2_0_COMB_FPDECODE_MOV5_1,
    I1 => GRLFPC2_0_COMB_FPDECODE_UN1_WREN210,
    I2 => GRLFPC2_0_COMB_FPDECODE_UN1_WREN210_1_0_0,
    I3 => GRLFPC2_0_MOV_2_SQMUXA_1_0,
    O => GRLFPC2_0_N_766);
  x_grlfpc2_0_comb_rs2_1_0x: LUT4 
  generic map(
    INIT => X"A0CC"
  )
  port map (
    I0 => cpi_d_inst(0),
    I1 => GRLFPC2_0_R_A_RS2(0),
    I2 => GRLFPC2_0_RS2_0_SQMUXA,
    I3 => holdn,
    O => GRLFPC2_0_COMB_RS2_1(0));
  x_grlfpc2_0_comb_rs2_1_1x: LUT4 
  generic map(
    INIT => X"A0CC"
  )
  port map (
    I0 => cpi_d_inst(1),
    I1 => GRLFPC2_0_R_A_RS2(1),
    I2 => GRLFPC2_0_RS2_0_SQMUXA,
    I3 => holdn,
    O => RFI2_RD2ADDR_0_INT_9_INT_21);
  x_grlfpc2_0_comb_rs2_1_2x: LUT4 
  generic map(
    INIT => X"A0CC"
  )
  port map (
    I0 => cpi_d_inst(2),
    I1 => GRLFPC2_0_R_A_RS2(2),
    I2 => GRLFPC2_0_RS2_0_SQMUXA,
    I3 => holdn,
    O => RFI2_RD2ADDR_1_INT_10_INT_22);
  x_grlfpc2_0_comb_rs2_1_3x: LUT4 
  generic map(
    INIT => X"A0CC"
  )
  port map (
    I0 => cpi_d_inst(3),
    I1 => GRLFPC2_0_R_A_RS2(3),
    I2 => GRLFPC2_0_RS2_0_SQMUXA,
    I3 => holdn,
    O => RFI2_RD2ADDR_2_INT_11_INT_23);
  x_grlfpc2_0_comb_rs2_1_4x: LUT4 
  generic map(
    INIT => X"A0CC"
  )
  port map (
    I0 => cpi_d_inst(4),
    I1 => GRLFPC2_0_R_A_RS2(4),
    I2 => GRLFPC2_0_RS2_0_SQMUXA,
    I3 => holdn,
    O => RFI2_RD2ADDR_3_INT_12_INT_24);
  x_grlfpc2_0_un1_afq6: LUT4 
  generic map(
    INIT => X"0E0F"
  )
  port map (
    I0 => cpi_d_inst(19),
    I1 => cpi_d_inst(20),
    I2 => GRLFPC2_0_AFQ_3_SQMUXA,
    I3 => GRLFPC2_0_COMB_FPDECODE_AFQ7_1,
    O => GRLFPC2_0_UN1_AFQ6_I);
  x_grlfpc2_0_comb_seqerr_un7_op: LUT2 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => GRLFPC2_0_COMB_SEQERR_UN13_OP,
    I1 => GRLFPC2_0_RS2_0_SQMUXA,
    O => GRLFPC2_0_COMB_SEQERR_UN7_OP_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_1_29x: LUT4 
  generic map(
    INIT => X"2000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTXZYFROMD_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(29),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_1(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_1_30x: LUT4 
  generic map(
    INIT => X"2000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTXZYFROMD_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(30),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_1(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_1_31x: LUT4 
  generic map(
    INIT => X"2000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTXZYFROMD_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(31),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_1(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_1_35x: LUT4 
  generic map(
    INIT => X"2000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTXZYFROMD_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(35),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_1(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_1_45x: LUT4 
  generic map(
    INIT => X"2000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTXZYFROMD_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(45),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_1(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_1_49x: LUT4 
  generic map(
    INIT => X"2000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTXZYFROMD_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(49),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_1(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_1_51x: LUT4 
  generic map(
    INIT => X"2000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTXZYFROMD_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_1(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_1_53x: LUT4 
  generic map(
    INIT => X"2000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTXZYFROMD_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_1(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_1_54x: LUT4 
  generic map(
    INIT => X"2000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTXZYFROMD_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(54),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_1(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_0_25x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP2(32),
    I2 => rfo2_data2(29),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_0_24x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP2(33),
    I2 => rfo2_data2(30),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_0_23x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP2(34),
    I2 => rfo2_data2(31),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_0_22x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP2(32),
    I2 => GRLFPC2_0_OP2(35),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_0_18x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP2(36),
    I2 => GRLFPC2_0_OP2(39),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_0_17x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP2(37),
    I2 => GRLFPC2_0_OP2(40),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_0_16x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP2(38),
    I2 => GRLFPC2_0_OP2(41),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_0_10x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP2(44),
    I2 => GRLFPC2_0_OP2(47),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_0_5x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP2(49),
    I2 => GRLFPC2_0_OP2(52),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_0_82x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP1(33),
    I2 => rfo2_data1(30),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(82));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_0_79x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP1(33),
    I2 => GRLFPC2_0_OP1(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(79));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_0_77x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP1(35),
    I2 => GRLFPC2_0_OP1(38),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(77));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_0_75x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP1(37),
    I2 => GRLFPC2_0_OP1(40),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(75));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_0_74x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP1(38),
    I2 => GRLFPC2_0_OP1(41),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(74));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_0_73x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP1(39),
    I2 => GRLFPC2_0_OP1(42),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(73));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_0_71x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP1(41),
    I2 => GRLFPC2_0_OP1(44),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(71));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_0_69x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP1(43),
    I2 => GRLFPC2_0_OP1(46),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(69));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_0_68x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP1(44),
    I2 => GRLFPC2_0_OP1(47),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(68));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_0_65x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP1(47),
    I2 => GRLFPC2_0_OP1(50),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(65));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_0_63x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP1(49),
    I2 => GRLFPC2_0_OP1(52),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(63));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_0_62x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP1(50),
    I2 => GRLFPC2_0_OP1(53),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(62));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_3x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_110,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(54),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_4x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_111,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_5x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_112,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(52),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_12x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_119,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(45),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_13x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_120,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(44),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_14x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_121,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(43),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_15x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_122,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(42),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_16x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_123,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(41),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_18x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_125,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(39),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_19x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_126,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(38),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_20x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_127,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(37),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_21x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_128,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(36),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_22x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_129,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(35),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_25x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_132,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(32),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_26x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_133,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(31),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_27x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_134,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(30),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_28x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_135,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(29),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_30x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_137,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(27),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_31x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_138,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(26),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_32x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_139,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(25),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_33x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_140,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(24),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_34x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_141,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_35x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_142,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(22),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_36x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_143,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_37x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_144,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(20),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_38x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_145,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_39x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_146,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(18),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_40x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_147,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_41x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_148,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(16),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_42x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_149,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(15),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_43x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_150,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(14),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_47x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_154,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(10),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_49x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_156,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_50x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_157,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(7),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_51x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_158,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(6),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_52x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_159,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_54x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_161,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_55x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_162,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(2),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_257x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I1 => GRLFPC2_0_OP1(52),
    I2 => GRLFPC2_0_OP1(55),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_377);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_256x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I1 => GRLFPC2_0_OP1(53),
    I2 => GRLFPC2_0_OP1(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_378);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_254x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I1 => GRLFPC2_0_OP1(55),
    I2 => GRLFPC2_0_OP1(58),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_380);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_253x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I1 => GRLFPC2_0_OP1(56),
    I2 => GRLFPC2_0_OP1(59),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_381);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_251x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I1 => GRLFPC2_0_OP1(58),
    I2 => GRLFPC2_0_OP1(61),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_383);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_250x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I1 => GRLFPC2_0_OP1(59),
    I2 => GRLFPC2_0_OP1(62),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_384);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_244x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(10),
    I2 => GRLFPC2_0_OP2(55),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_763);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_243x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(9),
    I2 => GRLFPC2_0_OP2(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_764);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_242x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
    I2 => GRLFPC2_0_OP2(57),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_765);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_241x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(7),
    I2 => GRLFPC2_0_OP2(58),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_766);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_239x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5),
    I2 => GRLFPC2_0_OP2(60),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_768);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_238x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
    I2 => GRLFPC2_0_OP2(61),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_769);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_237x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
    I2 => GRLFPC2_0_OP2(62),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_770);
  x_grlfpc2_0_wrdata_0_63x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(31),
    I1 => GRLFPC2_0_N_126,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_1_48x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_155,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(9),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_0_81x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP1(34),
    I2 => rfo2_data1(31),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(81));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_252x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I1 => GRLFPC2_0_OP1(57),
    I2 => GRLFPC2_0_OP1(60),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_382);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_255x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I1 => GRLFPC2_0_OP1(54),
    I2 => GRLFPC2_0_OP1(57),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_379);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_1_56x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_163,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_1_46x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_153,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(11),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_1_17x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_124,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(40),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_1_24x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_131,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(33),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_1_23x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_130,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(34),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_1_29x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_136,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(28),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_0_78x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP1(34),
    I2 => GRLFPC2_0_OP1(37),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(78));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_0_19x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP2(35),
    I2 => GRLFPC2_0_OP2(38),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_0_61x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP1(51),
    I2 => GRLFPC2_0_OP1(54),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(61));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_0_4x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP2(50),
    I2 => GRLFPC2_0_OP2(53),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_44x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_151,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(13),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_1_53x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_160,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_1_45x: LUT3_L 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_152,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(12),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_19_0_83x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP1(32),
    I2 => rfo2_data1(29),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(83));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_240x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(6),
    I2 => GRLFPC2_0_OP2(59),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_767);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_entryshft_un1_entrypoint: LUT4 
  generic map(
    INIT => X"0040"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN1_S_14,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(78),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(82),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(85),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN1_ENTRYPOINT);
  x_grlfpc2_0_comb_rsdecode_rs1v2: LUT2 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_FPDECODE_MOV5,
    I1 => GRLFPC2_0_COMB_RSDECODE_RS1V2_0,
    O => GRLFPC2_0_N_764);
  x_grlfpc2_0_mov_2_sqmuxa: LUT4 
  generic map(
    INIT => X"8000"
  )
  port map (
    I0 => GRLFPC2_0_COMB_FPDECODE_MOV11,
    I1 => GRLFPC2_0_MOV_2_SQMUXA_1_0,
    I2 => GRLFPC2_0_MOV_2_SQMUXA_1_1,
    I3 => GRLFPC2_0_MOV_2_SQMUXA_2,
    O => GRLFPC2_0_MOV_2_SQMUXA);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_un24_shdvar: LUT4 
  generic map(
    INIT => X"8000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(2),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(3),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN24_SHDVAR);
  x_grlfpc2_0_un1_afq7_i_a2_0: LUT4 
  generic map(
    INIT => X"8ACF"
  )
  port map (
    I0 => cpi_d_inst(6),
    I1 => cpi_d_inst(30),
    I2 => GRLFPC2_0_COMB_FPDECODE_MOV6,
    I3 => GRLFPC2_0_MOV_0_SQMUXA_2_0,
    O => GRLFPC2_0_UN1_AFQ7_I_A2_0);
  x_grlfpc2_0_un1_wren210_4_0: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_RS1V10_I,
    I1 => GRLFPC2_0_RS1V_1_SQMUXA,
    O => GRLFPC2_0_UN1_WREN210_4_0);
  x_grlfpc2_0_comb_v_i_v6_0: LUT4 
  generic map(
    INIT => X"CC08"
  )
  port map (
    I0 => GRLFPC2_0_R_I_EXEC,
    I1 => GRLFPC2_0_R_I_V,
    I2 => GRLFPC2_0_V_FSR_FTT_1_SQMUXA_2_2,
    I3 => GRLFPC2_0_V_I_EXEC_0_SQMUXA,
    O => GRLFPC2_0_COMB_V_I_V6_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_entryshft_entrypoint_2: LUT4 
  generic map(
    INIT => X"002A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_ENTRYPOINT_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN4_S_SQRT_1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN9_S_11_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN14_S_MOV,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_ENTRYPOINT_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_un7_shdvar: LUT4 
  generic map(
    INIT => X"00CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1870);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_117_1: LUT3 
  generic map(
    INIT => X"A6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_CIN_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(316),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2122_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_7: LUT4 
  generic map(
    INIT => X"6C93"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1019,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_8: LUT4 
  generic map(
    INIT => X"6C93"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1020,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_8);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_9: LUT4 
  generic map(
    INIT => X"6C93"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1021,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(9),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_9);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m14_0_1x: MUXF6 port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M13(1),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M12(1),
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SS12,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M14(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m14_0_2x: MUXF6 port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M13(2),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M12(2),
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SS12,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M14(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_57x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(174),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m14_0_0x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M12(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M13(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SS12,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M14(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_62_1_51x: LUT2 
  generic map(
    INIT => X"6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_CIN_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_114_1_1_0(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_62_1(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_98_1_0: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(29),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(344),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_98_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_108_0_5x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(12),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(361),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_50(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_64_0_49x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(56),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_CIN_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(317),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_6(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_107_0_6x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(13),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(360),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_49(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_101_0_12x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(19),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(354),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_43(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_61_1_0: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(43),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(330),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_61_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_88_1_0: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(32),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(341),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_88_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_62_1_0: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(28),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(345),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_62_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_94_0_19x: LUT3 
  generic map(
    INIT => X"96"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(26),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(26),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_36(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_89_0_24x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(31),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(342),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_31(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_97_0_16x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(350),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_39(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_85_0_28x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(35),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(338),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_27(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_90_0_23x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(343),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_32(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_74_1_0: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(38),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(335),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_74_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_81_0_32x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(39),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(334),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_23(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_86_0_27x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(34),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(339),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_28(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_74_0_39x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(46),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(327),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_16(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_96_1_0: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(48),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(325),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_96_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_76_0_37x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(44),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(329),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_18(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_78_0_35x: LUT3 
  generic map(
    INIT => X"96"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(42),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_20(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_83_0_30x: LUT3 
  generic map(
    INIT => X"96"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(37),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(37),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_25(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_104_0_9x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(16),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(357),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_46(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_75_0_38x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(45),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(328),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_17(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_95_0_18x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(25),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(348),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_37(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_87_0_26x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(33),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(340),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_29(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_64_1_0: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(52),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_CIN_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(321),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_64_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_si_113_0_0x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(7),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_CIN_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(366),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_113_0(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_SBLSBs_1_0_1x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(367),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SBLSBS_1_0(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_69_0_44x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(51),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(322),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_11(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_80_0_33x: LUT3 
  generic map(
    INIT => X"96"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(40),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_22(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_103_0_10x: LUT3 
  generic map(
    INIT => X"96"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(17),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_45(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_100_1_0: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(24),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_CIN_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(349),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_100_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_100_0_13x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(20),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(353),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_42(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_98_0_15x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(22),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_19_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(351),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_40(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_111_0_2x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(9),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_CIN_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(364),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_53(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_84_0_29x: LUT3 
  generic map(
    INIT => X"96"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(36),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(36),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_26(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_70_0_43x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(50),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(323),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_12(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_106_0_7x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(14),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_CIN_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(359),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_48(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_78_1_0: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(41),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(332),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_78_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_104_1_0: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(10),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(363),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_104_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_109_0_4x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(11),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_CIN_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(362),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_51(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_66_1_0: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(27),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(346),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_66_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_94_1_0: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(49),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(324),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_94_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_73_0_40x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(47),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(326),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_15(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_13_0: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(365),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_13_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_SBLSBs_0_0x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(5),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_CIN_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(368),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SBLSBS_0(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_67_0_46x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(53),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(320),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_9(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_65_0_48x: LUT3 
  generic map(
    INIT => X"96"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(55),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_7(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_105_0_8x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(15),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_CIN_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(358),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_47(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_66_0_47x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(54),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(319),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_8(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_102_0_11x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(18),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(355),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_44(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_99_0_14x: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_18_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(352),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_41(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_123: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_CIN_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(370),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SALSBS(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_114_0: LUT2 
  generic map(
    INIT => X"6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_CIN_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_114_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_1_0_4x: LUT2 
  generic map(
    INIT => X"6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_CIN_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_1_0(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_NE_2: LUT4_L 
  generic map(
    INIT => X"2112"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_5,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_1(6),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_NE_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_49_1_0_258x: LUT2_L 
  generic map(
    INIT => X"6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_CIN_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_114_1_1_0(56),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_49_1_0(258));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_m_6x: LUT4 
  generic map(
    INIT => X"5410"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I2 => GRLFPC2_0_OP2(48),
    I3 => GRLFPC2_0_OP2(51),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_m_3x: LUT4 
  generic map(
    INIT => X"5410"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I2 => GRLFPC2_0_OP2(51),
    I3 => GRLFPC2_0_OP2(54),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_m_9x: LUT4 
  generic map(
    INIT => X"5410"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I2 => GRLFPC2_0_OP2(45),
    I3 => GRLFPC2_0_OP2(48),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_m_20x: LUT4 
  generic map(
    INIT => X"5410"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I2 => GRLFPC2_0_OP2(34),
    I3 => GRLFPC2_0_OP2(37),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_1_0x: LUT4 
  generic map(
    INIT => X"6000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTXZYFROMD_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_m_7x: LUT4 
  generic map(
    INIT => X"5410"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I2 => GRLFPC2_0_OP2(47),
    I3 => GRLFPC2_0_OP2(50),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_v_1x: LUT4 
  generic map(
    INIT => X"738C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_2_1(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(56),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN20_XZXBUS(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_m_8x: LUT4 
  generic map(
    INIT => X"5410"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I2 => GRLFPC2_0_OP2(46),
    I3 => GRLFPC2_0_OP2(49),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_m_11x: LUT4 
  generic map(
    INIT => X"5410"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I2 => GRLFPC2_0_OP2(43),
    I3 => GRLFPC2_0_OP2(46),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_m_12x: LUT4 
  generic map(
    INIT => X"5410"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I2 => GRLFPC2_0_OP2(42),
    I3 => GRLFPC2_0_OP2(45),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_m_13x: LUT4 
  generic map(
    INIT => X"5410"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I2 => GRLFPC2_0_OP2(41),
    I3 => GRLFPC2_0_OP2(44),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_m_14x: LUT4 
  generic map(
    INIT => X"5410"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I2 => GRLFPC2_0_OP2(40),
    I3 => GRLFPC2_0_OP2(43),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_m_15x: LUT4 
  generic map(
    INIT => X"5410"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I2 => GRLFPC2_0_OP2(39),
    I3 => GRLFPC2_0_OP2(42),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_m_21x: LUT4 
  generic map(
    INIT => X"5410"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I2 => GRLFPC2_0_OP2(33),
    I3 => GRLFPC2_0_OP2(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M(21));
  x_grlfpc2_0_I_162_266: LUT4 
  generic map(
    INIT => X"00FE"
  )
  port map (
    I0 => N_2291_TZ,
    I1 => GRLFPC2_0_R_I_EXEC,
    I2 => GRLFPC2_0_R_X_FPOP,
    I3 => GRLFPC2_0_V_FSR_FTT_1_SQMUXA_2_2,
    O => GRLFPC2_0_N_791);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_7x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(7),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(11),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12120);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_7x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(9),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(13),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12121);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_7x: MUXF5 port map (
      I0 => N_12120,
      I1 => N_12121,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_8x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12122);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_8x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(10),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(14),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12123);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_8x: MUXF5 port map (
      I0 => N_12122,
      I1 => N_12123,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_9x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(9),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(13),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12124);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_9x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(11),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(15),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12125);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_9x: MUXF5 port map (
      I0 => N_12124,
      I1 => N_12125,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_10x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(10),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(14),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12126);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_10x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(12),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12127);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_10x: MUXF5 port map (
      I0 => N_12126,
      I1 => N_12127,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_11x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(11),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(13),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_12x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(12),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12128);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_12x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(14),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(18),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12129);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_12x: MUXF5 port map (
      I0 => N_12128,
      I1 => N_12129,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_13x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(13),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(15),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_14x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(14),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(18),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12130);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_14x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(16),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(20),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12131);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_14x: MUXF5 port map (
      I0 => N_12130,
      I1 => N_12131,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_15x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(15),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(17),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_16x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(16),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(20),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12132);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_16x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(18),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(22),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12133);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_16x: MUXF5 port map (
      I0 => N_12132,
      I1 => N_12133,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_18x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(18),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(22),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12134);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_18x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(20),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(24),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12135);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_18x: MUXF5 port map (
      I0 => N_12134,
      I1 => N_12135,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_19x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(19),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(21),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_20x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(20),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(22),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_21x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(21),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(23),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_22x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(22),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(24),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_23x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(27),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12136);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_23x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(25),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12137);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_23x: MUXF5 port map (
      I0 => N_12136,
      I1 => N_12137,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_24x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(24),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(26),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_25x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(25),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12138);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_25x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(27),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(31),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12139);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_25x: MUXF5 port map (
      I0 => N_12138,
      I1 => N_12139,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_26x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(26),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12140);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_26x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(28),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(32),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12141);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_26x: MUXF5 port map (
      I0 => N_12140,
      I1 => N_12141,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_27x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(27),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(31),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12142);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_27x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(29),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(33),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12143);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_27x: MUXF5 port map (
      I0 => N_12142,
      I1 => N_12143,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_28x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(28),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(32),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12144);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_28x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(34),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12145);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_28x: MUXF5 port map (
      I0 => N_12144,
      I1 => N_12145,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_29x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(29),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(33),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12146);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_29x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(31),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(35),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12147);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_29x: MUXF5 port map (
      I0 => N_12146,
      I1 => N_12147,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_30x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(34),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12148);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_30x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(32),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(36),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12149);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_30x: MUXF5 port map (
      I0 => N_12148,
      I1 => N_12149,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_31x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(31),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(35),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12150);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_31x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(33),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(37),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12151);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_31x: MUXF5 port map (
      I0 => N_12150,
      I1 => N_12151,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_32x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(32),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(36),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12152);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_32x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(34),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(38),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12153);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_32x: MUXF5 port map (
      I0 => N_12152,
      I1 => N_12153,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_33x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(33),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(37),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12154);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_33x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(35),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12155);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_33x: MUXF5 port map (
      I0 => N_12154,
      I1 => N_12155,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_34x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(34),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(38),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12156);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_34x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(36),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12157);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_34x: MUXF5 port map (
      I0 => N_12156,
      I1 => N_12157,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_40x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(42),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_42x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(44),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_46x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(46),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(48),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_48x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(48),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(52),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12158);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_48x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(50),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(54),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12159);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_48x: MUXF5 port map (
      I0 => N_12158,
      I1 => N_12159,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_49x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(49),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(51),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_50x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(50),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(54),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12160);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_50x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(52),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(56),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12161);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_50x: MUXF5 port map (
      I0 => N_12160,
      I1 => N_12161,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_51x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(53),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_52x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(52),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(56),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12162);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_52x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(54),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(57),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12163);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_52x: MUXF5 port map (
      I0 => N_12162,
      I1 => N_12163,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_53x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(55),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_54x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(54),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m14_0_bm_3x: LUT4 
  generic map(
    INIT => X"F7FF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SM0_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SM3_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV_4_0,
    O => N_12165);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m14_0_3x: MUXF5 port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M14_0X(3),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M14_0X_0(3),
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV_6,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M14(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_229x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_225);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_228x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(3),
    O => GRLFPC2_0_FPO_FRAC(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_227x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(4),
    O => GRLFPC2_0_FPO_FRAC(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_226x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(5),
    O => GRLFPC2_0_FPO_FRAC(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_225x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(6),
    O => GRLFPC2_0_FPO_FRAC(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_223x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(8),
    O => GRLFPC2_0_FPO_FRAC(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_222x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(9),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(9),
    O => GRLFPC2_0_FPO_FRAC(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_221x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(10),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(10),
    O => GRLFPC2_0_FPO_FRAC(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_220x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(11),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(11),
    O => GRLFPC2_0_FPO_FRAC(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_219x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(12),
    O => GRLFPC2_0_FPO_FRAC(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_218x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(13),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(13),
    O => GRLFPC2_0_FPO_FRAC(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_216x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(15),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(15),
    O => GRLFPC2_0_FPO_FRAC(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_215x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(16),
    O => GRLFPC2_0_FPO_FRAC(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_213x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(18),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(18),
    O => GRLFPC2_0_FPO_FRAC(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_212x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(19),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(19),
    O => GRLFPC2_0_FPO_FRAC(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_211x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(20),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(20),
    O => GRLFPC2_0_FPO_FRAC(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_210x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(21),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(21),
    O => GRLFPC2_0_FPO_FRAC(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_208x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(23),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(23),
    O => GRLFPC2_0_FPO_FRAC(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_205x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(26),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(26),
    O => GRLFPC2_0_FPO_FRAC(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_204x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(27),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(27),
    O => GRLFPC2_0_FPO_FRAC(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_203x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(28),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(28),
    O => GRLFPC2_0_FPO_FRAC(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_202x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(29),
    O => GRLFPC2_0_FPO_FRAC(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_201x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(30),
    O => GRLFPC2_0_FPO_FRAC(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_200x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(31),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(31),
    O => GRLFPC2_0_FPO_FRAC(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_199x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(32),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(32),
    O => GRLFPC2_0_FPO_FRAC(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_198x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(33),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(33),
    O => GRLFPC2_0_FPO_FRAC(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_197x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(34),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(34),
    O => GRLFPC2_0_FPO_FRAC(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_196x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(35),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(35),
    O => GRLFPC2_0_FPO_FRAC(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_195x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(36),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(36),
    O => GRLFPC2_0_FPO_FRAC(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_192x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(39),
    O => GRLFPC2_0_FPO_FRAC(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_191x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(40),
    O => GRLFPC2_0_FPO_FRAC(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_190x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(41),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(41),
    O => GRLFPC2_0_FPO_FRAC(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_189x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(42),
    O => GRLFPC2_0_FPO_FRAC(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_188x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(43),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(43),
    O => GRLFPC2_0_FPO_FRAC(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_187x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(44),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(44),
    O => GRLFPC2_0_FPO_FRAC(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_186x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(45),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(45),
    O => GRLFPC2_0_FPO_FRAC(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_185x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(46),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(46),
    O => GRLFPC2_0_FPO_FRAC(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_179x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(52),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(52),
    O => GRLFPC2_0_FPO_FRAC(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_175x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(56),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_279);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_i_m2_0_224x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(7),
    O => GRLFPC2_0_FPO_FRAC(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_i_m2_0_209x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(22),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(22),
    O => GRLFPC2_0_FPO_FRAC(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_i_m2_0_207x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(24),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(24),
    O => GRLFPC2_0_FPO_FRAC(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_t_3_i_m2_0_0x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(57),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(57),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2276);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_i_m2_0_184x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(47),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(47),
    O => GRLFPC2_0_FPO_FRAC(47));
  x_grlfpc2_0_comb_v_i_res_1_0_am_52x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_EXP(0),
    I2 => GRLFPC2_0_R_I_RES(52),
    O => N_12166);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_52x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(23),
    I2 => rfo2_data2(23),
    O => N_12167);
  x_grlfpc2_0_comb_v_i_res_1_0_52x: MUXF5 port map (
      I0 => N_12166,
      I1 => N_12167,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(52));
  x_grlfpc2_0_comb_v_i_res_1_0_am_53x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_EXP(1),
    I2 => GRLFPC2_0_R_I_RES(53),
    O => N_12168);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_53x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(24),
    I2 => rfo2_data2(24),
    O => N_12169);
  x_grlfpc2_0_comb_v_i_res_1_0_53x: MUXF5 port map (
      I0 => N_12168,
      I1 => N_12169,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(53));
  x_grlfpc2_0_comb_v_i_res_1_0_am_54x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_EXP(2),
    I2 => GRLFPC2_0_R_I_RES(54),
    O => N_12170);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_54x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(25),
    I2 => rfo2_data2(25),
    O => N_12171);
  x_grlfpc2_0_comb_v_i_res_1_0_54x: MUXF5 port map (
      I0 => N_12170,
      I1 => N_12171,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(54));
  x_grlfpc2_0_comb_v_i_res_1_0_am_55x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_EXP(3),
    I2 => GRLFPC2_0_R_I_RES(55),
    O => N_12172);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_55x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(26),
    I2 => rfo2_data2(26),
    O => N_12173);
  x_grlfpc2_0_comb_v_i_res_1_0_55x: MUXF5 port map (
      I0 => N_12172,
      I1 => N_12173,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(55));
  x_grlfpc2_0_comb_v_i_res_1_0_am_56x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_EXP(4),
    I2 => GRLFPC2_0_R_I_RES(56),
    O => N_12174);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_56x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(27),
    I2 => rfo2_data2(27),
    O => N_12175);
  x_grlfpc2_0_comb_v_i_res_1_0_56x: MUXF5 port map (
      I0 => N_12174,
      I1 => N_12175,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(56));
  x_grlfpc2_0_comb_v_i_res_1_0_am_57x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_EXP(5),
    I2 => GRLFPC2_0_R_I_RES(57),
    O => N_12176);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_57x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(28),
    I2 => rfo2_data2(28),
    O => N_12177);
  x_grlfpc2_0_comb_v_i_res_1_0_57x: MUXF5 port map (
      I0 => N_12176,
      I1 => N_12177,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(57));
  x_grlfpc2_0_comb_v_i_res_1_0_am_58x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_EXP(6),
    I2 => GRLFPC2_0_R_I_RES(58),
    O => N_12178);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_58x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(29),
    I2 => rfo2_data2(29),
    O => N_12179);
  x_grlfpc2_0_comb_v_i_res_1_0_58x: MUXF5 port map (
      I0 => N_12178,
      I1 => N_12179,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(58));
  x_grlfpc2_0_comb_v_i_res_1_0_am_59x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_EXP(7),
    I2 => GRLFPC2_0_R_I_RES(59),
    O => N_12180);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_59x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(30),
    I2 => rfo2_data2(30),
    O => N_12181);
  x_grlfpc2_0_comb_v_i_res_1_0_59x: MUXF5 port map (
      I0 => N_12180,
      I1 => N_12181,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(59));
  x_grlfpc2_0_comb_wrdata_4_0_0x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(0),
    I2 => GRLFPC2_0_R_I_RES(29),
    O => GRLFPC2_0_COMB_WRDATA_4(0));
  x_grlfpc2_0_comb_wrdata_4_0_2x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(2),
    I2 => GRLFPC2_0_R_I_RES(31),
    O => GRLFPC2_0_COMB_WRDATA_4(2));
  x_grlfpc2_0_comb_wrdata_4_0_4x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(4),
    I2 => GRLFPC2_0_R_I_RES(33),
    O => GRLFPC2_0_COMB_WRDATA_4(4));
  x_grlfpc2_0_comb_wrdata_4_0_5x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(5),
    I2 => GRLFPC2_0_R_I_RES(34),
    O => GRLFPC2_0_COMB_WRDATA_4(5));
  x_grlfpc2_0_comb_wrdata_4_0_6x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(6),
    I2 => GRLFPC2_0_R_I_RES(35),
    O => GRLFPC2_0_COMB_WRDATA_4(6));
  x_grlfpc2_0_comb_wrdata_4_0_7x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(7),
    I2 => GRLFPC2_0_R_I_RES(36),
    O => GRLFPC2_0_COMB_WRDATA_4(7));
  x_grlfpc2_0_comb_wrdata_4_0_8x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(8),
    I2 => GRLFPC2_0_R_I_RES(37),
    O => GRLFPC2_0_COMB_WRDATA_4(8));
  x_grlfpc2_0_comb_wrdata_4_0_9x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(9),
    I2 => GRLFPC2_0_R_I_RES(38),
    O => GRLFPC2_0_COMB_WRDATA_4(9));
  x_grlfpc2_0_comb_wrdata_4_0_10x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(10),
    I2 => GRLFPC2_0_R_I_RES(39),
    O => GRLFPC2_0_COMB_WRDATA_4(10));
  x_grlfpc2_0_comb_wrdata_4_0_11x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(11),
    I2 => GRLFPC2_0_R_I_RES(40),
    O => GRLFPC2_0_COMB_WRDATA_4(11));
  x_grlfpc2_0_comb_wrdata_4_0_12x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(12),
    I2 => GRLFPC2_0_R_I_RES(41),
    O => GRLFPC2_0_COMB_WRDATA_4(12));
  x_grlfpc2_0_comb_wrdata_4_0_14x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(14),
    I2 => GRLFPC2_0_R_I_RES(43),
    O => GRLFPC2_0_COMB_WRDATA_4(14));
  x_grlfpc2_0_comb_wrdata_4_0_15x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(15),
    I2 => GRLFPC2_0_R_I_RES(44),
    O => GRLFPC2_0_COMB_WRDATA_4(15));
  x_grlfpc2_0_comb_wrdata_4_0_18x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(18),
    I2 => GRLFPC2_0_R_I_RES(47),
    O => GRLFPC2_0_COMB_WRDATA_4(18));
  x_grlfpc2_0_comb_wrdata_4_0_19x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(19),
    I2 => GRLFPC2_0_R_I_RES(48),
    O => GRLFPC2_0_COMB_WRDATA_4(19));
  x_grlfpc2_0_comb_wrdata_4_0_21x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(21),
    I2 => GRLFPC2_0_R_I_RES(50),
    O => GRLFPC2_0_COMB_WRDATA_4(21));
  x_grlfpc2_0_comb_wrdata_4_0_22x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(22),
    I2 => GRLFPC2_0_R_I_RES(51),
    O => GRLFPC2_0_COMB_WRDATA_4(22));
  x_grlfpc2_0_comb_wrdata_4_0_23x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(23),
    I2 => GRLFPC2_0_R_I_RES(52),
    O => GRLFPC2_0_COMB_WRDATA_4(23));
  x_grlfpc2_0_comb_wrdata_4_0_24x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(24),
    I2 => GRLFPC2_0_R_I_RES(53),
    O => GRLFPC2_0_COMB_WRDATA_4(24));
  x_grlfpc2_0_comb_wrdata_4_0_25x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(25),
    I2 => GRLFPC2_0_R_I_RES(54),
    O => GRLFPC2_0_COMB_WRDATA_4(25));
  x_grlfpc2_0_comb_wrdata_4_0_26x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(26),
    I2 => GRLFPC2_0_R_I_RES(55),
    O => GRLFPC2_0_COMB_WRDATA_4(26));
  x_grlfpc2_0_comb_wrdata_4_0_28x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(28),
    I2 => GRLFPC2_0_R_I_RES(57),
    O => GRLFPC2_0_COMB_WRDATA_4(28));
  x_grlfpc2_0_comb_wrdata_4_0_29x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(29),
    I2 => GRLFPC2_0_R_I_RES(58),
    O => GRLFPC2_0_COMB_WRDATA_4(29));
  x_grlfpc2_0_comb_wrdata_4_0_31x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(31),
    I2 => GRLFPC2_0_R_I_RES(63),
    O => GRLFPC2_0_COMB_WRDATA_4(31));
  x_grlfpc2_0_comb_wrdata_4_0_32x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(29),
    I2 => GRLFPC2_0_R_I_RES(32),
    O => GRLFPC2_0_COMB_WRDATA_4(32));
  x_grlfpc2_0_comb_wrdata_4_0_34x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(31),
    I2 => GRLFPC2_0_R_I_RES(34),
    O => GRLFPC2_0_COMB_WRDATA_4(34));
  x_grlfpc2_0_comb_wrdata_4_0_36x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(33),
    I2 => GRLFPC2_0_R_I_RES(36),
    O => GRLFPC2_0_COMB_WRDATA_4(36));
  x_grlfpc2_0_comb_wrdata_4_0_37x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(34),
    I2 => GRLFPC2_0_R_I_RES(37),
    O => GRLFPC2_0_COMB_WRDATA_4(37));
  x_grlfpc2_0_comb_wrdata_4_0_38x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(35),
    I2 => GRLFPC2_0_R_I_RES(38),
    O => GRLFPC2_0_COMB_WRDATA_4(38));
  x_grlfpc2_0_comb_wrdata_4_0_39x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(36),
    I2 => GRLFPC2_0_R_I_RES(39),
    O => GRLFPC2_0_COMB_WRDATA_4(39));
  x_grlfpc2_0_comb_wrdata_4_0_40x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(37),
    I2 => GRLFPC2_0_R_I_RES(40),
    O => GRLFPC2_0_COMB_WRDATA_4(40));
  x_grlfpc2_0_comb_wrdata_4_0_41x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(38),
    I2 => GRLFPC2_0_R_I_RES(41),
    O => GRLFPC2_0_COMB_WRDATA_4(41));
  x_grlfpc2_0_comb_wrdata_4_0_42x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(39),
    I2 => GRLFPC2_0_R_I_RES(42),
    O => GRLFPC2_0_COMB_WRDATA_4(42));
  x_grlfpc2_0_comb_wrdata_4_0_43x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(40),
    I2 => GRLFPC2_0_R_I_RES(43),
    O => GRLFPC2_0_COMB_WRDATA_4(43));
  x_grlfpc2_0_comb_wrdata_4_0_44x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(41),
    I2 => GRLFPC2_0_R_I_RES(44),
    O => GRLFPC2_0_COMB_WRDATA_4(44));
  x_grlfpc2_0_comb_wrdata_4_0_46x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(43),
    I2 => GRLFPC2_0_R_I_RES(46),
    O => GRLFPC2_0_COMB_WRDATA_4(46));
  x_grlfpc2_0_comb_wrdata_4_0_47x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(44),
    I2 => GRLFPC2_0_R_I_RES(47),
    O => GRLFPC2_0_COMB_WRDATA_4(47));
  x_grlfpc2_0_comb_wrdata_4_0_50x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(47),
    I2 => GRLFPC2_0_R_I_RES(50),
    O => GRLFPC2_0_COMB_WRDATA_4(50));
  x_grlfpc2_0_comb_wrdata_4_0_51x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(48),
    I2 => GRLFPC2_0_R_I_RES(51),
    O => GRLFPC2_0_COMB_WRDATA_4(51));
  x_grlfpc2_0_comb_wrdata_4_0_53x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(50),
    I2 => GRLFPC2_0_R_I_RES(53),
    O => GRLFPC2_0_COMB_WRDATA_4(53));
  x_grlfpc2_0_comb_wrdata_4_0_54x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(51),
    I2 => GRLFPC2_0_R_I_RES(54),
    O => GRLFPC2_0_COMB_WRDATA_4(54));
  x_grlfpc2_0_comb_wrdata_4_0_55x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(52),
    I2 => GRLFPC2_0_R_I_RES(55),
    O => GRLFPC2_0_COMB_WRDATA_4(55));
  x_grlfpc2_0_comb_wrdata_4_0_56x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(53),
    I2 => GRLFPC2_0_R_I_RES(56),
    O => GRLFPC2_0_COMB_WRDATA_4(56));
  x_grlfpc2_0_comb_wrdata_4_0_57x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(54),
    I2 => GRLFPC2_0_R_I_RES(57),
    O => GRLFPC2_0_COMB_WRDATA_4(57));
  x_grlfpc2_0_comb_wrdata_4_0_58x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(55),
    I2 => GRLFPC2_0_R_I_RES(58),
    O => GRLFPC2_0_COMB_WRDATA_4(58));
  x_grlfpc2_0_comb_wrdata_4_0_60x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(57),
    I2 => GRLFPC2_0_R_I_RES(60),
    O => GRLFPC2_0_COMB_WRDATA_4(60));
  x_grlfpc2_0_comb_wrdata_4_0_61x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(58),
    I2 => GRLFPC2_0_R_I_RES(61),
    O => GRLFPC2_0_COMB_WRDATA_4(61));
  x_grlfpc2_0_wraddr_1_0_1x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_addr(1),
    I1 => GRLFPC2_0_COMB_WRADDR_5(1),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => RFI2_WRADDR_0_INT_13_INT_25);
  x_grlfpc2_0_wraddr_1_0_2x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_addr(2),
    I1 => GRLFPC2_0_COMB_WRADDR_5(2),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => RFI2_WRADDR_1_INT_14_INT_26);
  x_grlfpc2_0_wraddr_1_0_3x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_addr(3),
    I1 => GRLFPC2_0_COMB_WRADDR_5(3),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => RFI2_WRADDR_2_INT_15_INT_27);
  x_grlfpc2_0_wraddr_1_0_4x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_addr(4),
    I1 => GRLFPC2_0_COMB_WRADDR_5(4),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => RFI2_WRADDR_3_INT_16_INT_28);
  x_grlfpc2_0_comb_v_e_stdata_1_0_am_12x: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(44),
    I1 => GRLFPC2_0_R_A_AFSR,
    O => N_12182);
  x_grlfpc2_0_comb_v_e_stdata_1_0_bm_12x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(12),
    I2 => GRLFPC2_0_R_I_PC(12),
    O => N_12183);
  x_grlfpc2_0_comb_v_e_stdata_1_0_12x: MUXF5 port map (
      I0 => N_12182,
      I1 => N_12183,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(12));
  x_grlfpc2_0_comb_v_e_stdata_1_0_am_15x: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(47),
    I1 => GRLFPC2_0_R_A_AFSR,
    O => N_12184);
  x_grlfpc2_0_comb_v_e_stdata_1_0_bm_15x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(15),
    I2 => GRLFPC2_0_R_I_PC(15),
    O => N_12185);
  x_grlfpc2_0_comb_v_e_stdata_1_0_15x: MUXF5 port map (
      I0 => N_12184,
      I1 => N_12185,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(15));
  x_grlfpc2_0_comb_v_e_stdata_1_0_am_17x: LUT2 
  generic map(
    INIT => X"E"
  )
  port map (
    I0 => GRLFPC2_0_OP1(49),
    I1 => GRLFPC2_0_R_A_AFSR,
    O => N_12186);
  x_grlfpc2_0_comb_v_e_stdata_1_0_bm_17x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(17),
    I2 => GRLFPC2_0_R_I_PC(17),
    O => N_12187);
  x_grlfpc2_0_comb_v_e_stdata_1_0_17x: MUXF5 port map (
      I0 => N_12186,
      I1 => N_12187,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(17));
  x_grlfpc2_0_comb_v_e_stdata_1_0_am_18x: LUT2 
  generic map(
    INIT => X"E"
  )
  port map (
    I0 => GRLFPC2_0_OP1(50),
    I1 => GRLFPC2_0_R_A_AFSR,
    O => N_12188);
  x_grlfpc2_0_comb_v_e_stdata_1_0_bm_18x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(18),
    I2 => GRLFPC2_0_R_I_PC(18),
    O => N_12189);
  x_grlfpc2_0_comb_v_e_stdata_1_0_18x: MUXF5 port map (
      I0 => N_12188,
      I1 => N_12189,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(18));
  x_grlfpc2_0_comb_v_e_stdata_1_0_am_21x: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(53),
    I1 => GRLFPC2_0_R_A_AFSR,
    O => N_12190);
  x_grlfpc2_0_comb_v_e_stdata_1_0_bm_21x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(21),
    I2 => GRLFPC2_0_R_I_PC(21),
    O => N_12191);
  x_grlfpc2_0_comb_v_e_stdata_1_0_21x: MUXF5 port map (
      I0 => N_12190,
      I1 => N_12191,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(21));
  x_grlfpc2_0_comb_v_e_stdata_1_0_am_29x: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(61),
    I1 => GRLFPC2_0_R_A_AFSR,
    O => N_12192);
  x_grlfpc2_0_comb_v_e_stdata_1_0_bm_29x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(29),
    I2 => GRLFPC2_0_R_I_PC(29),
    O => N_12193);
  x_grlfpc2_0_comb_v_e_stdata_1_0_29x: MUXF5 port map (
      I0 => N_12192,
      I1 => N_12193,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_181x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(50),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(50),
    O => GRLFPC2_0_FPO_FRAC(50));
  x_grlfpc2_0_comb_wrdata_4_0_62x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(59),
    I2 => GRLFPC2_0_R_I_RES(62),
    O => GRLFPC2_0_COMB_WRDATA_4(62));
  x_grlfpc2_0_comb_wrdata_4_0_59x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(56),
    I2 => GRLFPC2_0_R_I_RES(59),
    O => GRLFPC2_0_COMB_WRDATA_4(59));
  x_grlfpc2_0_comb_wrdata_4_0_33x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(30),
    I2 => GRLFPC2_0_R_I_RES(33),
    O => GRLFPC2_0_COMB_WRDATA_4(33));
  x_grlfpc2_0_comb_wrdata_4_0_30x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(30),
    I2 => GRLFPC2_0_R_I_RES(59),
    O => GRLFPC2_0_COMB_WRDATA_4(30));
  x_grlfpc2_0_comb_wrdata_4_0_27x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(27),
    I2 => GRLFPC2_0_R_I_RES(56),
    O => GRLFPC2_0_COMB_WRDATA_4(27));
  x_grlfpc2_0_comb_wrdata_4_0_1x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(1),
    I2 => GRLFPC2_0_R_I_RES(30),
    O => GRLFPC2_0_COMB_WRDATA_4(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_i_m2_0_182x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(49),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(49),
    O => GRLFPC2_0_FPO_FRAC(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_230x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_224);
  x_grlfpc2_0_comb_v_e_stdata_1_2_am_28x: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(60),
    I1 => GRLFPC2_0_R_A_AFSR,
    O => N_12194);
  x_grlfpc2_0_comb_v_e_stdata_1_2_bm_28x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(28),
    I2 => GRLFPC2_0_R_I_PC(28),
    O => N_12195);
  x_grlfpc2_0_comb_v_e_stdata_1_2_28x: MUXF5 port map (
      I0 => N_12194,
      I1 => N_12195,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_231x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_223);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_1x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12196);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_1x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12197);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_1x: MUXF5 port map (
      I0 => N_12196,
      I1 => N_12197,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_0x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12198);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_0x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12199);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_0x: MUXF5 port map (
      I0 => N_12198,
      I1 => N_12199,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_217x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(14),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(14),
    O => GRLFPC2_0_FPO_FRAC(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_35x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(35),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12200);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_35x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(37),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(41),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12201);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_35x: MUXF5 port map (
      I0 => N_12200,
      I1 => N_12201,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_5x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(5),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(9),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12202);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_5x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(7),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(11),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12203);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_5x: MUXF5 port map (
      I0 => N_12202,
      I1 => N_12203,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_4x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(4),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12204);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_4x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(10),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12205);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_4x: MUXF5 port map (
      I0 => N_12204,
      I1 => N_12205,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_3x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12206);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_3x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(5),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(9),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12207);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_3x: MUXF5 port map (
      I0 => N_12206,
      I1 => N_12207,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_2x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12208);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_2x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(4),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12209);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_2x: MUXF5 port map (
      I0 => N_12208,
      I1 => N_12209,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_214x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(17),
    O => GRLFPC2_0_FPO_FRAC(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_i_m2_0_206x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(25),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(25),
    O => GRLFPC2_0_FPO_FRAC(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_194x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(37),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(37),
    O => GRLFPC2_0_FPO_FRAC(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_193x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(38),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(38),
    O => GRLFPC2_0_FPO_FRAC(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_17x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(19),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_183x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(48),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(48),
    O => GRLFPC2_0_FPO_FRAC(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_38x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(38),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12210);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_38x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(40),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(44),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12211);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_38x: MUXF5 port map (
      I0 => N_12210,
      I1 => N_12211,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_36x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(36),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(38),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_i_m2_0_180x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(51),
    O => GRLFPC2_0_FPO_FRAC(51));
  x_grlfpc2_0_comb_v_e_stdata_1_0_am_19x: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(51),
    I1 => GRLFPC2_0_R_A_AFSR,
    O => N_12212);
  x_grlfpc2_0_comb_v_e_stdata_1_0_bm_19x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(19),
    I2 => GRLFPC2_0_R_I_PC(19),
    O => N_12213);
  x_grlfpc2_0_comb_v_e_stdata_1_0_19x: MUXF5 port map (
      I0 => N_12212,
      I1 => N_12213,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(19));
  x_grlfpc2_0_comb_v_e_stdata_1_2_am_20x: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(52),
    I1 => GRLFPC2_0_R_A_AFSR,
    O => N_12214);
  x_grlfpc2_0_comb_v_e_stdata_1_2_bm_20x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(20),
    I2 => GRLFPC2_0_R_I_PC(20),
    O => N_12215);
  x_grlfpc2_0_comb_v_e_stdata_1_2_20x: MUXF5 port map (
      I0 => N_12214,
      I1 => N_12215,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_i_m2_0_178x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(53),
    O => GRLFPC2_0_FPO_FRAC(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_43x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(43),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(45),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_177x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(54),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(54),
    O => GRLFPC2_0_FPO_FRAC(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_am_47x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(47),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12216);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_bm_47x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(49),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12217);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_47x: MUXF5 port map (
      I0 => N_12216,
      I1 => N_12217,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_45x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(45),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(47),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_41x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(41),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(43),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_37x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(37),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(39),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(37));
  x_grlfpc2_0_comb_wrdata_4_0_52x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(49),
    I2 => GRLFPC2_0_R_I_RES(52),
    O => GRLFPC2_0_COMB_WRDATA_4(52));
  x_grlfpc2_0_comb_wrdata_4_0_49x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(46),
    I2 => GRLFPC2_0_R_I_RES(49),
    O => GRLFPC2_0_COMB_WRDATA_4(49));
  x_grlfpc2_0_comb_wrdata_4_0_48x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(45),
    I2 => GRLFPC2_0_R_I_RES(48),
    O => GRLFPC2_0_COMB_WRDATA_4(48));
  x_grlfpc2_0_comb_wrdata_4_0_45x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(42),
    I2 => GRLFPC2_0_R_I_RES(45),
    O => GRLFPC2_0_COMB_WRDATA_4(45));
  x_grlfpc2_0_comb_wrdata_4_0_35x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(32),
    I2 => GRLFPC2_0_R_I_RES(35),
    O => GRLFPC2_0_COMB_WRDATA_4(35));
  x_grlfpc2_0_comb_wrdata_4_0_20x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(20),
    I2 => GRLFPC2_0_R_I_RES(49),
    O => GRLFPC2_0_COMB_WRDATA_4(20));
  x_grlfpc2_0_comb_wrdata_4_0_17x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(17),
    I2 => GRLFPC2_0_R_I_RES(46),
    O => GRLFPC2_0_COMB_WRDATA_4(17));
  x_grlfpc2_0_comb_wrdata_4_0_16x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(16),
    I2 => GRLFPC2_0_R_I_RES(45),
    O => GRLFPC2_0_COMB_WRDATA_4(16));
  x_grlfpc2_0_comb_wrdata_4_0_13x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(13),
    I2 => GRLFPC2_0_R_I_RES(42),
    O => GRLFPC2_0_COMB_WRDATA_4(13));
  x_grlfpc2_0_comb_wrdata_4_0_3x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_R_I_RES(3),
    I2 => GRLFPC2_0_R_I_RES(32),
    O => GRLFPC2_0_COMB_WRDATA_4(3));
  x_grlfpc2_0_comb_v_i_v6: LUT4 
  generic map(
    INIT => X"EF00"
  )
  port map (
    I0 => GRLFPC2_0_COMB_MEXC_1(0),
    I1 => GRLFPC2_0_COMB_MEXC_1(1),
    I2 => GRLFPC2_0_COMB_UN1_MEXC_2,
    I3 => GRLFPC2_0_COMB_V_I_V6_0,
    O => GRLFPC2_0_COMB_V_I_V6);
  x_grlfpc2_0_comb_wren2_9_iv_0: LUT4 
  generic map(
    INIT => X"45CF"
  )
  port map (
    I0 => cpi_x_inst(25),
    I1 => GRLFPC2_0_COMB_WREN22,
    I2 => GRLFPC2_0_WREN2_1_SQMUXA_1_0,
    I3 => GRLFPC2_0_WREN2_2_SQMUXA,
    O => GRLFPC2_0_COMB_WREN2_9_IV_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_21x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(36),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(210),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_45x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(12),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(186),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_6x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(225),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_46x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(11),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(185),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_5x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(52),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(226),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_14x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(43),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(217),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_2x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(229),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_20x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(37),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(211),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_53x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(178),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_25x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(32),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(206),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_56x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(175),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_15x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(42),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(216),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_44x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(13),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(187),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_13x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(44),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(218),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_7x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(50),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(224),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_8x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(49),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(223),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_19x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(38),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(212),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_51x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(6),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(180),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_49x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(182),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_55x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(2),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(176),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_38x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(193),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_35x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(22),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(196),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_29x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(28),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(202),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_52x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(179),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_50x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(7),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(181),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_12x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(45),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(219),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_31x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(26),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(200),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_17x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(40),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(214),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_42x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(15),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(189),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_47x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(10),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(184),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_10x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(47),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(221),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_3x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(54),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(228),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_40x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(191),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_18x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(39),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(213),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_37x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(20),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(194),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_16x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(41),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(215),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_23x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(34),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(208),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_39x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(18),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(192),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_30x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(27),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(201),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_11x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(46),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(220),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_54x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(177),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_22x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(35),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(209),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_27x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(30),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(204),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_4x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(227),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_24x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(33),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(207),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_36x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(195),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_48x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(9),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(183),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_34x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(197),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_43x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(14),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(188),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_41x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(16),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(190),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_9x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(48),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(222),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_33x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(24),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(198),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_32x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(25),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(199),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_26x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(31),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(205),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_0_28x: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS25,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS26,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(29),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(203),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(28));
  x_grlfpc2_0_comb_v_e_stdata_1_1_am_0x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(32),
    I1 => GRLFPC2_0_R_A_AFSR,
    I2 => GRLFPC2_0_R_FSR_CEXC(0),
    O => N_12218);
  x_grlfpc2_0_comb_v_e_stdata_1_1_0x: MUXF5 port map (
      I0 => N_12218,
      I1 => N_12219,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(0));
  x_grlfpc2_0_comb_v_e_stdata_1_0_am_2x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(34),
    I1 => GRLFPC2_0_R_A_AFSR,
    I2 => GRLFPC2_0_R_FSR_CEXC(2),
    O => N_12220);
  x_grlfpc2_0_comb_v_e_stdata_1_0_bm_2x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(2),
    I2 => GRLFPC2_0_R_I_PC(2),
    O => N_12221);
  x_grlfpc2_0_comb_v_e_stdata_1_0_2x: MUXF5 port map (
      I0 => N_12220,
      I1 => N_12221,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(2));
  x_grlfpc2_0_comb_v_e_stdata_1_0_am_3x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(35),
    I1 => GRLFPC2_0_R_A_AFSR,
    I2 => GRLFPC2_0_R_FSR_CEXC(3),
    O => N_12222);
  x_grlfpc2_0_comb_v_e_stdata_1_0_bm_3x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(3),
    I2 => GRLFPC2_0_R_I_PC(3),
    O => N_12223);
  x_grlfpc2_0_comb_v_e_stdata_1_0_3x: MUXF5 port map (
      I0 => N_12222,
      I1 => N_12223,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(3));
  x_grlfpc2_0_comb_v_e_stdata_1_0_am_4x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(36),
    I1 => GRLFPC2_0_R_A_AFSR,
    I2 => GRLFPC2_0_R_FSR_CEXC(4),
    O => N_12224);
  x_grlfpc2_0_comb_v_e_stdata_1_0_bm_4x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(4),
    I2 => GRLFPC2_0_R_I_PC(4),
    O => N_12225);
  x_grlfpc2_0_comb_v_e_stdata_1_0_4x: MUXF5 port map (
      I0 => N_12224,
      I1 => N_12225,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(4));
  x_grlfpc2_0_comb_v_e_stdata_1_0_am_5x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(37),
    I1 => GRLFPC2_0_R_A_AFSR,
    I2 => GRLFPC2_0_R_FSR_AEXC(0),
    O => N_12226);
  x_grlfpc2_0_comb_v_e_stdata_1_0_bm_5x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(5),
    I2 => GRLFPC2_0_R_I_PC(5),
    O => N_12227);
  x_grlfpc2_0_comb_v_e_stdata_1_0_5x: MUXF5 port map (
      I0 => N_12226,
      I1 => N_12227,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(5));
  x_grlfpc2_0_comb_v_e_stdata_1_0_am_6x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(38),
    I1 => GRLFPC2_0_R_A_AFSR,
    I2 => GRLFPC2_0_R_FSR_AEXC(1),
    O => N_12228);
  x_grlfpc2_0_comb_v_e_stdata_1_0_bm_6x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(6),
    I2 => GRLFPC2_0_R_I_PC(6),
    O => N_12229);
  x_grlfpc2_0_comb_v_e_stdata_1_0_6x: MUXF5 port map (
      I0 => N_12228,
      I1 => N_12229,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(6));
  x_grlfpc2_0_comb_v_e_stdata_1_0_am_7x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(39),
    I1 => GRLFPC2_0_R_A_AFSR,
    I2 => GRLFPC2_0_R_FSR_AEXC(2),
    O => N_12230);
  x_grlfpc2_0_comb_v_e_stdata_1_0_bm_7x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(7),
    I2 => GRLFPC2_0_R_I_PC(7),
    O => N_12231);
  x_grlfpc2_0_comb_v_e_stdata_1_0_7x: MUXF5 port map (
      I0 => N_12230,
      I1 => N_12231,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(7));
  x_grlfpc2_0_comb_v_e_stdata_1_0_am_8x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(40),
    I1 => GRLFPC2_0_R_A_AFSR,
    I2 => GRLFPC2_0_R_FSR_AEXC(3),
    O => N_12232);
  x_grlfpc2_0_comb_v_e_stdata_1_0_bm_8x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(8),
    I2 => GRLFPC2_0_R_I_PC(8),
    O => N_12233);
  x_grlfpc2_0_comb_v_e_stdata_1_0_8x: MUXF5 port map (
      I0 => N_12232,
      I1 => N_12233,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(8));
  x_grlfpc2_0_comb_v_e_stdata_1_0_am_9x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(41),
    I1 => GRLFPC2_0_R_A_AFSR,
    I2 => GRLFPC2_0_R_FSR_AEXC(4),
    O => N_12234);
  x_grlfpc2_0_comb_v_e_stdata_1_0_bm_9x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(9),
    I2 => GRLFPC2_0_R_I_PC(9),
    O => N_12235);
  x_grlfpc2_0_comb_v_e_stdata_1_0_9x: MUXF5 port map (
      I0 => N_12234,
      I1 => N_12235,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(9));
  x_grlfpc2_0_comb_v_e_stdata_1_0_am_10x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => CPO_CC_0_INT_3,
    I1 => GRLFPC2_0_OP1(42),
    I2 => GRLFPC2_0_R_A_AFSR,
    O => N_12236);
  x_grlfpc2_0_comb_v_e_stdata_1_0_bm_10x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(10),
    I2 => GRLFPC2_0_R_I_PC(10),
    O => N_12237);
  x_grlfpc2_0_comb_v_e_stdata_1_0_10x: MUXF5 port map (
      I0 => N_12236,
      I1 => N_12237,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(10));
  x_grlfpc2_0_comb_v_e_stdata_1_0_am_11x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => CPO_CC_1_INT_4,
    I1 => GRLFPC2_0_OP1(43),
    I2 => GRLFPC2_0_R_A_AFSR,
    O => N_12238);
  x_grlfpc2_0_comb_v_e_stdata_1_0_bm_11x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(11),
    I2 => GRLFPC2_0_R_I_PC(11),
    O => N_12239);
  x_grlfpc2_0_comb_v_e_stdata_1_0_11x: MUXF5 port map (
      I0 => N_12238,
      I1 => N_12239,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(11));
  x_grlfpc2_0_comb_v_e_stdata_1_0_am_13x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(45),
    I1 => GRLFPC2_0_R_A_AFSR,
    I2 => GRLFPC2_0_SEQERR_1_SQMUXA_1_SN,
    O => N_12240);
  x_grlfpc2_0_comb_v_e_stdata_1_0_bm_13x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(13),
    I2 => GRLFPC2_0_R_I_PC(13),
    O => N_12241);
  x_grlfpc2_0_comb_v_e_stdata_1_0_13x: MUXF5 port map (
      I0 => N_12240,
      I1 => N_12241,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(13));
  x_grlfpc2_0_comb_v_e_stdata_1_0_am_14x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(46),
    I1 => GRLFPC2_0_R_A_AFSR,
    I2 => GRLFPC2_0_R_FSR_FTT(0),
    O => N_12242);
  x_grlfpc2_0_comb_v_e_stdata_1_0_bm_14x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(14),
    I2 => GRLFPC2_0_R_I_PC(14),
    O => N_12243);
  x_grlfpc2_0_comb_v_e_stdata_1_0_14x: MUXF5 port map (
      I0 => N_12242,
      I1 => N_12243,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(14));
  x_grlfpc2_0_comb_v_e_stdata_1_0_am_16x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(48),
    I1 => GRLFPC2_0_R_A_AFSR,
    I2 => GRLFPC2_0_R_FSR_FTT(2),
    O => N_12244);
  x_grlfpc2_0_comb_v_e_stdata_1_0_bm_16x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(16),
    I2 => GRLFPC2_0_R_I_PC(16),
    O => N_12245);
  x_grlfpc2_0_comb_v_e_stdata_1_0_16x: MUXF5 port map (
      I0 => N_12244,
      I1 => N_12245,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(16));
  x_grlfpc2_0_comb_v_e_stdata_1_0_am_23x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(55),
    I1 => GRLFPC2_0_R_A_AFSR,
    I2 => GRLFPC2_0_R_FSR_TEM(0),
    O => N_12246);
  x_grlfpc2_0_comb_v_e_stdata_1_0_bm_23x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(23),
    I2 => GRLFPC2_0_R_I_PC(23),
    O => N_12247);
  x_grlfpc2_0_comb_v_e_stdata_1_0_23x: MUXF5 port map (
      I0 => N_12246,
      I1 => N_12247,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(23));
  x_grlfpc2_0_comb_v_e_stdata_1_0_am_27x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(59),
    I1 => GRLFPC2_0_R_A_AFSR,
    I2 => GRLFPC2_0_R_FSR_TEM(4),
    O => N_12248);
  x_grlfpc2_0_comb_v_e_stdata_1_0_bm_27x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(27),
    I2 => GRLFPC2_0_R_I_PC(27),
    O => N_12249);
  x_grlfpc2_0_comb_v_e_stdata_1_0_27x: MUXF5 port map (
      I0 => N_12248,
      I1 => N_12249,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(27));
  x_grlfpc2_0_comb_v_e_stdata_1_0_am_31x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(63),
    I1 => GRLFPC2_0_R_A_AFSR,
    I2 => GRLFPC2_0_R_FSR_RD(1),
    O => N_12250);
  x_grlfpc2_0_comb_v_e_stdata_1_0_bm_31x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(31),
    I2 => GRLFPC2_0_R_I_PC(31),
    O => N_12251);
  x_grlfpc2_0_comb_v_e_stdata_1_0_31x: MUXF5 port map (
      I0 => N_12250,
      I1 => N_12251,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(31));
  x_grlfpc2_0_comb_v_e_stdata_1_2_am_26x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(58),
    I1 => GRLFPC2_0_R_A_AFSR,
    I2 => GRLFPC2_0_R_FSR_TEM(3),
    O => N_12252);
  x_grlfpc2_0_comb_v_e_stdata_1_2_bm_26x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(26),
    I2 => GRLFPC2_0_R_I_PC(26),
    O => N_12253);
  x_grlfpc2_0_comb_v_e_stdata_1_2_26x: MUXF5 port map (
      I0 => N_12252,
      I1 => N_12253,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(26));
  x_grlfpc2_0_comb_v_e_stdata_1_0_am_25x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(57),
    I1 => GRLFPC2_0_R_A_AFSR,
    I2 => GRLFPC2_0_R_FSR_TEM(2),
    O => N_12254);
  x_grlfpc2_0_comb_v_e_stdata_1_0_bm_25x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(25),
    I2 => GRLFPC2_0_R_I_PC(25),
    O => N_12255);
  x_grlfpc2_0_comb_v_e_stdata_1_0_25x: MUXF5 port map (
      I0 => N_12254,
      I1 => N_12255,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(25));
  x_grlfpc2_0_comb_v_e_stdata_1_2_am_1x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(33),
    I1 => GRLFPC2_0_R_A_AFSR,
    I2 => GRLFPC2_0_R_FSR_CEXC(1),
    O => N_12256);
  x_grlfpc2_0_comb_v_e_stdata_1_2_1x: MUXF5 port map (
      I0 => N_12256,
      I1 => N_12257,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(1));
  x_grlfpc2_0_comb_rs1d_1_m2_0_0: LUT4 
  generic map(
    INIT => X"ACAA"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RS1D_1_M1,
    I1 => GRLFPC2_0_MOV_3_SQMUXA_1,
    I2 => GRLFPC2_0_MOV_7_SQMUXA,
    I3 => GRLFPC2_0_UN1_AFQ3_I,
    O => GRLFPC2_0_COMB_RS1D_1_M2);
  x_grlfpc2_0_I_231_0: LUT3 
  generic map(
    INIT => X"8B"
  )
  port map (
    I0 => cpi_d_inst(25),
    I1 => cpi_d_inst(30),
    I2 => GRLFPC2_0_N_764,
    O => GRLFPC2_0_N_674);
  x_grlfpc2_0_comb_v_e_stdata_1_2_am_22x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(54),
    I1 => GRLFPC2_0_R_A_AFSR,
    I2 => GRLFPC2_0_R_FSR_NONSTD,
    O => N_12258);
  x_grlfpc2_0_comb_v_e_stdata_1_2_bm_22x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(22),
    I2 => GRLFPC2_0_R_I_PC(22),
    O => N_12259);
  x_grlfpc2_0_comb_v_e_stdata_1_2_22x: MUXF5 port map (
      I0 => N_12258,
      I1 => N_12259,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(22));
  x_grlfpc2_0_comb_v_e_stdata_1_2_am_30x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(62),
    I1 => GRLFPC2_0_R_A_AFSR,
    I2 => GRLFPC2_0_R_FSR_RD(0),
    O => N_12260);
  x_grlfpc2_0_comb_v_e_stdata_1_2_bm_30x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(30),
    I2 => GRLFPC2_0_R_I_PC(30),
    O => N_12261);
  x_grlfpc2_0_comb_v_e_stdata_1_2_30x: MUXF5 port map (
      I0 => N_12260,
      I1 => N_12261,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(30));
  x_grlfpc2_0_comb_v_e_stdata_1_2_am_24x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_OP1(56),
    I1 => GRLFPC2_0_R_A_AFSR,
    I2 => GRLFPC2_0_R_FSR_TEM(1),
    O => N_12262);
  x_grlfpc2_0_comb_v_e_stdata_1_2_bm_24x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_E_STDATA2,
    I1 => GRLFPC2_0_R_I_INST(24),
    I2 => GRLFPC2_0_R_I_PC(24),
    O => N_12263);
  x_grlfpc2_0_comb_v_e_stdata_1_2_24x: MUXF5 port map (
      I0 => N_12262,
      I1 => N_12263,
      S => GRLFPC2_0_R_A_AFQ,
      O => GRLFPC2_0_COMB_V_E_STDATA_1(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_temp_1_1_1x: LUT4 
  generic map(
    INIT => X"00E0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_CIN_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(370),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => N_8928);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_13: LUT2 
  generic map(
    INIT => X"6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_13_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_15);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_waitmulxff_notsampledwait: LUT4 
  generic map(
    INIT => X"C808"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN17_WQSTSETS,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT);
  x_grlfpc2_0_I_223: LUT3 
  generic map(
    INIT => X"01"
  )
  port map (
    I0 => cpi_d_inst(14),
    I1 => cpi_d_inst(30),
    I2 => GRLFPC2_0_N_673,
    O => GRLFPC2_0_N_670);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_121_0_0_48x: LUT3 
  generic map(
    INIT => X"96"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_CIN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_114_1_1_0(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_121_0(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_NE_4: LUT4 
  generic map(
    INIT => X"8000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_11_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_12_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_NE_0,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_NE_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_NE_4);
  x_grlfpc2_0_v_state_2_sqmuxa: LUT3 
  generic map(
    INIT => X"31"
  )
  port map (
    I0 => GRLFPC2_0_N_781,
    I1 => GRLFPC2_0_COMB_V_I_V6,
    I2 => GRLFPC2_0_V_STATE_1_SQMUXA_1,
    O => GRLFPC2_0_V_STATE_2_SQMUXA);
  x_grlfpc2_0_comb_un1_r_i_v_1_264: LUT4 
  generic map(
    INIT => X"5504"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_I_V6,
    I1 => GRLFPC2_0_R_I_EXEC,
    I2 => GRLFPC2_0_V_FSR_FTT_1_SQMUXA_2_2,
    I3 => GRLFPC2_0_V_I_EXEC_0_SQMUXA,
    O => GRLFPC2_0_N_789);
  x_grlfpc2_0_v_fsr_ftt_1_sqmuxa_2_1: LUT2_L 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_I_V6,
    I1 => rst,
    LO => GRLFPC2_0_V_FSR_FTT_1_SQMUXA_2_1);
  x_grlfpc2_0_comb_seqerr_seqerrs2: LUT3 
  generic map(
    INIT => X"C5"
  )
  port map (
    I0 => GRLFPC2_0_AFQ_3_SQMUXA,
    I1 => GRLFPC2_0_COMB_SEQERR_UN7_OP_I,
    I2 => GRLFPC2_0_SEQERR_1_SQMUXA_1_SN,
    O => GRLFPC2_0_N_736);
  x_grlfpc2_0_comb_annulres_1_iv: LUT4 
  generic map(
    INIT => X"C8CC"
  )
  port map (
    I0 => GRLFPC2_0_N_781,
    I1 => GRLFPC2_0_N_791,
    I2 => GRLFPC2_0_R_I_EXEC,
    I3 => GRLFPC2_0_R_X_FPOP,
    O => GRLFPC2_0_V_I_EXEC26);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_0: LUT4_L 
  generic map(
    INIT => X"9C63"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN39_XZYBUSLSBS,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_2_1(0),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_0);
  x_grlfpc2_0_comb_v_i_res_1_0_am_63x: LUT3 
  generic map(
    INIT => X"72"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2000,
    I2 => GRLFPC2_0_R_I_RES(63),
    O => N_12264);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_63x: LUT3 
  generic map(
    INIT => X"12"
  )
  port map (
    I0 => cpi_a_inst(7),
    I1 => cpi_a_inst(8),
    I2 => GRLFPC2_0_OP2(63),
    O => N_12265);
  x_grlfpc2_0_comb_v_i_res_1_0_63x: MUXF5 port map (
      I0 => N_12264,
      I1 => N_12265,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(63));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_40x: LUT3_L 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(16),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1549);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_39x: LUT3_L 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1550);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_38x: LUT3_L 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(38),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(18),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1551);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_37x: LUT3_L 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(37),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1552);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_43x: LUT3_L 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(43),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(13),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1546);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_42x: LUT3 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(14),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1547);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_41x: LUT3_L 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(41),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(15),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1548);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_47x: LUT3_L 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(47),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(9),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1542);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_46x: LUT3_L 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(46),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(10),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1543);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_45x: LUT3_L 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(45),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(11),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1544);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_44x: LUT3 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(44),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(12),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1545);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_50x: LUT3_L 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(50),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(6),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1539);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_52x: LUT3_L 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(52),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1537);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_18x: LUT3 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(18),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(38),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1571);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_23x: LUT3 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(23),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(33),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1566);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_22x: LUT3 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(22),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(34),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1567);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_28x: LUT3 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(28),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(28),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1561);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_32x: LUT3_L 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(32),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(24),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1557);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_30x: LUT3 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(26),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1559);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_29x: LUT3 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(27),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1560);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_36x: LUT3_L 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(36),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(20),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1553);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_35x: LUT3_L 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(35),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1554);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_34x: LUT3_L 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(34),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(22),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1555);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_33x: LUT3_L 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(33),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1556);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_10x: LUT3 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(10),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(46),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1579);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_9x: LUT3 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(9),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(47),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1580);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_8x: LUT3 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(48),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1581);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_13x: LUT3 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(13),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(43),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1576);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_12x: LUT3 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(44),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1577);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_16x: LUT3 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(40),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1573);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_14x: LUT3 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(14),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(42),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1575);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_20x: LUT3 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(20),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1569);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_19x: LUT3 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(19),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(37),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1570);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_6x: LUT3 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(50),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1583);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_4x: LUT3 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(52),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1585);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_startshft_un3_notdecodedunimp: LUT4 
  generic map(
    INIT => X"0D00"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_ENTRYPOINT_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN1_ENTRYPOINT,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(65),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(67),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTDECODEDUNIMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_pctrl_new_14_77x: LUT4 
  generic map(
    INIT => X"2A00"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CONDMUXMULXFF_UN4_NOTSQRTLFTCC,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_OPREXCSHFT_UN3_OPREXC,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN42_CONDITIONAL,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(46),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14(77));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_56x: LUT3_L 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(56),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1533);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_54x: LUT3_L 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(54),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(2),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1535);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_55x: LUT3 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1534);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_48x: LUT3_L 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(48),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1541);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_49x: LUT3_L 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(49),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(7),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1540);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_51x: LUT3_L 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1538);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_iv_24x: LUT3 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(24),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(32),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1565);
  x_grlfpc2_0_un1_afq7_i_a2_2: LUT3 
  generic map(
    INIT => X"10"
  )
  port map (
    I0 => GRLFPC2_0_COMB_FPDECODE_AFQ7,
    I1 => GRLFPC2_0_MOV_3_SQMUXA_1,
    I2 => GRLFPC2_0_UN1_AFQ7_I_A2_0,
    O => GRLFPC2_0_UN1_AFQ7_I_A2_2);
  x_grlfpc2_0_comb_rdd_1_0_0: LUT4 
  generic map(
    INIT => X"2000"
  )
  port map (
    I0 => cpi_d_inst(31),
    I1 => GRLFPC2_0_RS1V_1_SQMUXA,
    I2 => GRLFPC2_0_UN1_AFQ3_I,
    I3 => GRLFPC2_0_UN1_AFQ6_I,
    O => GRLFPC2_0_COMB_RDD_1_0_0);
  x_grlfpc2_0_comb_v_a_afsr_1_0_1: LUT3 
  generic map(
    INIT => X"40"
  )
  port map (
    I0 => GRLFPC2_0_N_716,
    I1 => GRLFPC2_0_RS1V10_I,
    I2 => GRLFPC2_0_UN1_AFQ6_I,
    O => GRLFPC2_0_COMB_V_A_AFSR_1_0_1);
  x_grlfpc2_0_I_162_1: LUT3 
  generic map(
    INIT => X"40"
  )
  port map (
    I0 => GRLFPC2_0_N_691,
    I1 => GRLFPC2_0_N_791,
    I2 => rst,
    O => GRLFPC2_0_I_162_1);
  x_grlfpc2_0_comb_rs1d_1_0: LUT4 
  generic map(
    INIT => X"C0C8"
  )
  port map (
    I0 => cpi_d_inst(31),
    I1 => GRLFPC2_0_COMB_RS1D_1_M2,
    I2 => GRLFPC2_0_MOV_7_SQMUXA,
    I3 => GRLFPC2_0_RS1V_1_SQMUXA,
    O => GRLFPC2_0_COMB_RS1D_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_update_1: LUT2 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_pxs_multiplexormulxff_result_0_sn_m1_0_a3: LUT3 
  generic map(
    INIT => X"0D"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN1_MIFROMINST_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_71);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_52_CA_5_52x: LUT3 
  generic map(
    INIT => X"17"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(55),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1935);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_38_CA_19_38x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(41),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(332),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1949);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_39_CA_18_39x: LUT3 
  generic map(
    INIT => X"17"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(42),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1948);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_42_CA_15_42x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(45),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(328),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1945);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_45_CA_12_45x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(48),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(325),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1942);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_47_CA_10_47x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(50),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(323),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1940);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_48_CA_9_48x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(51),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(322),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1939);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_22_CA_35_22x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(25),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(348),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1965);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_CA_34_23x: LUT3 
  generic map(
    INIT => X"17"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(26),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(26),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1964);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_CA_33_24x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(27),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(346),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1963);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_25_CA_32_25x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(28),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(345),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1962);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_27_CA_30_27x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(343),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1960);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_28_CA_29_28x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(31),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(342),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1959);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_30_CA_27_30x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(33),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(340),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1957);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_31_CA_26_31x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(34),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(339),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1956);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_32_CA_25_32x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(35),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(338),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1955);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_34_CA_23_34x: LUT3 
  generic map(
    INIT => X"17"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(37),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(37),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1953);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_35_CA_22_35x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(38),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(335),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1952);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_CA_50_7x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(10),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(363),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1980);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_CA_47_10x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(13),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(360),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1977);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_CA_53_4x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(7),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_CIN_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(366),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1983);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_5_CA_52_5x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(365),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1982);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_53_CA_4_53x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(56),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_CIN_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(317),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1934);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_29_CA_28_29x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(32),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(341),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1958);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_CA_48_9x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(12),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(361),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1978);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_8_CA_49_8x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(11),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_CIN_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(362),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1979);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_6_CA_51_6x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(9),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_CIN_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(364),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1981);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_1_CA_56_1x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(4),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(369),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1987);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_20_CA_37_20x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(350),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1967);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_21_CA_36_21x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(24),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_CIN_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(349),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1966);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_44_CA_13_44x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(47),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(326),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1943);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_43_CA_14_43x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(46),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(327),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1944);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_37_CA_20_37x: LUT3 
  generic map(
    INIT => X"17"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(40),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1950);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_36_CA_21_36x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(39),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(334),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1951);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_33_CA_24_33x: LUT3 
  generic map(
    INIT => X"17"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(36),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(36),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1954);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_51_CA_6_51x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(54),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(319),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1936);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_50_CA_7_50x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(53),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(320),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1937);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_26_CA_31_26x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(29),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(344),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1961);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_14_CA_43_14x: LUT3 
  generic map(
    INIT => X"17"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(17),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1973);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_13_CA_44_13x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(16),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(357),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1974);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_49_CA_8_49x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(52),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_CIN_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(321),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1938);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_46_CA_11_46x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(49),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(324),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1941);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_19_CA_38_19x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(22),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_19_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(351),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1968);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_18_CA_39_18x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_18_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(352),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1969);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_17_CA_40_17x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(20),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(353),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1970);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_16_CA_41_16x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(19),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(354),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1971);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_15_CA_42_15x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(18),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(355),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1972);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_CA_54_3x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(367),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1984);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_CA_55_2x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(5),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_CIN_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(368),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1985);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_12_CA_45_12x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(15),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_CIN_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(358),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1975);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_CA_46_11x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(14),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_CIN_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(359),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1976);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_40_CA_17_40x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(43),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(330),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1947);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_41_CA_16_41x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(44),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(329),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1946);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notrembit_0_0x: LUT3 
  generic map(
    INIT => X"1D"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(52),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELINITREMBIT,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notrembit_0_1x: LUT3 
  generic map(
    INIT => X"1D"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(53),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELINITREMBIT,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notrembit_0_2x: LUT3 
  generic map(
    INIT => X"1D"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(54),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELINITREMBIT,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_notrembit_0_3x: LUT3 
  generic map(
    INIT => X"1D"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_278,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELINITREMBIT,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_1x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_2x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(3),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_3x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_5x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(6),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_6x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_7x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(8),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_8x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(9),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_9x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(9),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(10),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_10x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(10),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(11),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_11x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(11),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(12),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_12x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(13),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_13x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(13),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(14),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_14x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(14),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(15),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_17x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(18),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_18x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(18),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(19),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_19x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(19),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(20),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_20x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(20),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(21),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_21x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(21),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(22),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_22x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(22),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(23),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_23x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(23),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(24),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_24x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(24),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(25),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_25x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(25),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(26),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_26x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(26),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(27),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_27x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(27),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(28),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_28x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(28),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(29),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_29x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(30),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_30x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(31),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_31x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(31),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(32),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_32x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(32),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(33),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_33x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(33),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(34),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_34x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(34),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(35),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_35x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(35),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_36x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(36),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(37),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_37x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(37),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(38),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_am_38x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(38),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(40),
    O => N_12266);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_bm_38x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(41),
    O => N_12267);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_38x: MUXF5 port map (
      I0 => N_12266,
      I1 => N_12267,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_am_39x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(41),
    O => N_12268);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_bm_39x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(42),
    O => N_12269);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_39x: MUXF5 port map (
      I0 => N_12268,
      I1 => N_12269,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_40x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(41),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_41x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(41),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(42),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_42x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(43),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_am_43x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(43),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(45),
    O => N_12270);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_bm_43x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(44),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(46),
    O => N_12271);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_43x: MUXF5 port map (
      I0 => N_12270,
      I1 => N_12271,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_48x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(48),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(49),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_49x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(49),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(50),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_50x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(50),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(51),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_51x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(52),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_am_55x: LUT4 
  generic map(
    INIT => X"3335"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(55),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(57),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12272);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_bm_55x: LUT4 
  generic map(
    INIT => X"3335"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(56),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(57),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    O => N_12273);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_55x: MUXF5 port map (
      I0 => N_12272,
      I1 => N_12273,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_56x: LUT4 
  generic map(
    INIT => X"5754"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(57),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_17_0_0: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_279,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2276,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(52),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_363);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_112x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_224,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_566);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_110x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(3),
    I1 => GRLFPC2_0_FPO_FRAC(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_568);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_109x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(4),
    I1 => GRLFPC2_0_FPO_FRAC(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_569);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_108x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(5),
    I1 => GRLFPC2_0_FPO_FRAC(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_570);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_107x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(6),
    I1 => GRLFPC2_0_FPO_FRAC(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_571);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_105x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(8),
    I1 => GRLFPC2_0_FPO_FRAC(10),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_573);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_104x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(9),
    I1 => GRLFPC2_0_FPO_FRAC(11),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_574);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_103x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(10),
    I1 => GRLFPC2_0_FPO_FRAC(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_575);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_102x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(11),
    I1 => GRLFPC2_0_FPO_FRAC(13),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_576);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_101x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(12),
    I1 => GRLFPC2_0_FPO_FRAC(14),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_577);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_93x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(20),
    I1 => GRLFPC2_0_FPO_FRAC(22),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_585);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_92x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(21),
    I1 => GRLFPC2_0_FPO_FRAC(23),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_586);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_90x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(23),
    I1 => GRLFPC2_0_FPO_FRAC(25),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_588);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_88x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(25),
    I1 => GRLFPC2_0_FPO_FRAC(27),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_590);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_82x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(31),
    I1 => GRLFPC2_0_FPO_FRAC(33),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_596);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_79x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(34),
    I1 => GRLFPC2_0_FPO_FRAC(36),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_599);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_77x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(36),
    I1 => GRLFPC2_0_FPO_FRAC(38),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_601);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_75x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(38),
    I1 => GRLFPC2_0_FPO_FRAC(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_603);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_74x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(39),
    I1 => GRLFPC2_0_FPO_FRAC(41),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_604);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_73x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(40),
    I1 => GRLFPC2_0_FPO_FRAC(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_605);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_71x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(42),
    I1 => GRLFPC2_0_FPO_FRAC(44),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_607);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_69x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(44),
    I1 => GRLFPC2_0_FPO_FRAC(46),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_609);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_68x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(45),
    I1 => GRLFPC2_0_FPO_FRAC(47),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_610);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_63x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(50),
    I1 => GRLFPC2_0_FPO_FRAC(52),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_615);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_62x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(51),
    I1 => GRLFPC2_0_FPO_FRAC(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_616);
  x_grlfpc2_0_comb_v_i_res_3_0_32x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_FRAC(35),
    I2 => GRLFPC2_0_R_I_RES(32),
    LO => GRLFPC2_0_COMB_V_I_RES_3(32));
  x_grlfpc2_0_comb_v_i_res_3_0_33x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_FRAC(36),
    I2 => GRLFPC2_0_R_I_RES(33),
    LO => GRLFPC2_0_COMB_V_I_RES_3(33));
  x_grlfpc2_0_comb_v_i_res_3_0_35x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_FRAC(38),
    I2 => GRLFPC2_0_R_I_RES(35),
    LO => GRLFPC2_0_COMB_V_I_RES_3(35));
  x_grlfpc2_0_wrdata_0_0_0x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(0),
    I1 => GRLFPC2_0_COMB_WRDATA_4(0),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_63);
  x_grlfpc2_0_wrdata_0_0_2x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(2),
    I1 => GRLFPC2_0_COMB_WRDATA_4(2),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_65);
  x_grlfpc2_0_wrdata_0_0_4x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(4),
    I1 => GRLFPC2_0_COMB_WRDATA_4(4),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_67);
  x_grlfpc2_0_wrdata_0_0_5x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(5),
    I1 => GRLFPC2_0_COMB_WRDATA_4(5),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_68);
  x_grlfpc2_0_wrdata_0_0_6x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(6),
    I1 => GRLFPC2_0_COMB_WRDATA_4(6),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_69);
  x_grlfpc2_0_wrdata_0_0_7x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(7),
    I1 => GRLFPC2_0_COMB_WRDATA_4(7),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_70);
  x_grlfpc2_0_wrdata_0_0_8x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(8),
    I1 => GRLFPC2_0_COMB_WRDATA_4(8),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_71);
  x_grlfpc2_0_wrdata_0_0_9x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(9),
    I1 => GRLFPC2_0_COMB_WRDATA_4(9),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_72);
  x_grlfpc2_0_wrdata_0_0_10x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(10),
    I1 => GRLFPC2_0_COMB_WRDATA_4(10),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_73);
  x_grlfpc2_0_wrdata_0_0_11x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(11),
    I1 => GRLFPC2_0_COMB_WRDATA_4(11),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_74);
  x_grlfpc2_0_wrdata_0_0_12x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(12),
    I1 => GRLFPC2_0_COMB_WRDATA_4(12),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_75);
  x_grlfpc2_0_wrdata_0_0_14x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(14),
    I1 => GRLFPC2_0_COMB_WRDATA_4(14),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_77);
  x_grlfpc2_0_wrdata_0_0_15x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(15),
    I1 => GRLFPC2_0_COMB_WRDATA_4(15),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_78);
  x_grlfpc2_0_wrdata_0_0_18x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(18),
    I1 => GRLFPC2_0_COMB_WRDATA_4(18),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_81);
  x_grlfpc2_0_wrdata_0_0_19x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(19),
    I1 => GRLFPC2_0_COMB_WRDATA_4(19),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_82);
  x_grlfpc2_0_wrdata_0_0_21x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(21),
    I1 => GRLFPC2_0_COMB_WRDATA_4(21),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_84);
  x_grlfpc2_0_wrdata_0_0_22x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(22),
    I1 => GRLFPC2_0_COMB_WRDATA_4(22),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_85);
  x_grlfpc2_0_wrdata_0_0_23x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(23),
    I1 => GRLFPC2_0_COMB_WRDATA_4(23),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_86);
  x_grlfpc2_0_wrdata_0_0_24x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(24),
    I1 => GRLFPC2_0_COMB_WRDATA_4(24),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_87);
  x_grlfpc2_0_wrdata_0_0_25x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(25),
    I1 => GRLFPC2_0_COMB_WRDATA_4(25),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_88);
  x_grlfpc2_0_wrdata_0_0_26x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(26),
    I1 => GRLFPC2_0_COMB_WRDATA_4(26),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_89);
  x_grlfpc2_0_wrdata_0_0_28x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(28),
    I1 => GRLFPC2_0_COMB_WRDATA_4(28),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_91);
  x_grlfpc2_0_wrdata_0_0_29x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(29),
    I1 => GRLFPC2_0_COMB_WRDATA_4(29),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_92);
  x_grlfpc2_0_wrdata_0_0_31x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(31),
    I1 => GRLFPC2_0_COMB_WRDATA_4(31),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_94);
  x_grlfpc2_0_wrdata_0_0_32x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(0),
    I1 => GRLFPC2_0_COMB_WRDATA_4(32),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_95);
  x_grlfpc2_0_wrdata_0_0_34x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(2),
    I1 => GRLFPC2_0_COMB_WRDATA_4(34),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_97);
  x_grlfpc2_0_wrdata_0_0_36x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(4),
    I1 => GRLFPC2_0_COMB_WRDATA_4(36),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_99);
  x_grlfpc2_0_wrdata_0_0_37x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(5),
    I1 => GRLFPC2_0_COMB_WRDATA_4(37),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_100);
  x_grlfpc2_0_wrdata_0_0_38x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(6),
    I1 => GRLFPC2_0_COMB_WRDATA_4(38),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_101);
  x_grlfpc2_0_wrdata_0_0_39x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(7),
    I1 => GRLFPC2_0_COMB_WRDATA_4(39),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_102);
  x_grlfpc2_0_wrdata_0_0_40x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(8),
    I1 => GRLFPC2_0_COMB_WRDATA_4(40),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_103);
  x_grlfpc2_0_wrdata_0_0_41x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(9),
    I1 => GRLFPC2_0_COMB_WRDATA_4(41),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_104);
  x_grlfpc2_0_wrdata_0_0_42x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(10),
    I1 => GRLFPC2_0_COMB_WRDATA_4(42),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_105);
  x_grlfpc2_0_wrdata_0_0_43x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(11),
    I1 => GRLFPC2_0_COMB_WRDATA_4(43),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_106);
  x_grlfpc2_0_wrdata_0_0_44x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(12),
    I1 => GRLFPC2_0_COMB_WRDATA_4(44),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_107);
  x_grlfpc2_0_wrdata_0_0_46x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(14),
    I1 => GRLFPC2_0_COMB_WRDATA_4(46),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_109);
  x_grlfpc2_0_wrdata_0_0_47x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(15),
    I1 => GRLFPC2_0_COMB_WRDATA_4(47),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_110);
  x_grlfpc2_0_wrdata_0_0_50x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(18),
    I1 => GRLFPC2_0_COMB_WRDATA_4(50),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_113);
  x_grlfpc2_0_wrdata_0_0_51x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(19),
    I1 => GRLFPC2_0_COMB_WRDATA_4(51),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_114);
  x_grlfpc2_0_wrdata_0_0_53x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(21),
    I1 => GRLFPC2_0_COMB_WRDATA_4(53),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_116);
  x_grlfpc2_0_wrdata_0_0_54x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(22),
    I1 => GRLFPC2_0_COMB_WRDATA_4(54),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_117);
  x_grlfpc2_0_wrdata_0_0_55x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(23),
    I1 => GRLFPC2_0_COMB_WRDATA_4(55),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_118);
  x_grlfpc2_0_wrdata_0_0_56x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(24),
    I1 => GRLFPC2_0_COMB_WRDATA_4(56),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_119);
  x_grlfpc2_0_wrdata_0_0_57x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(25),
    I1 => GRLFPC2_0_COMB_WRDATA_4(57),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_120);
  x_grlfpc2_0_wrdata_0_0_58x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(26),
    I1 => GRLFPC2_0_COMB_WRDATA_4(58),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_121);
  x_grlfpc2_0_wrdata_0_0_60x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(28),
    I1 => GRLFPC2_0_COMB_WRDATA_4(60),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_123);
  x_grlfpc2_0_wrdata_0_0_61x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(29),
    I1 => GRLFPC2_0_COMB_WRDATA_4(61),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_124);
  x_grlfpc2_0_wrdata_0_0_62x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(30),
    I1 => GRLFPC2_0_COMB_WRDATA_4(62),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_125);
  x_grlfpc2_0_wrdata_0_0_59x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(27),
    I1 => GRLFPC2_0_COMB_WRDATA_4(59),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_122);
  x_grlfpc2_0_wrdata_0_0_33x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(1),
    I1 => GRLFPC2_0_COMB_WRDATA_4(33),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_96);
  x_grlfpc2_0_wrdata_0_0_30x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(30),
    I1 => GRLFPC2_0_COMB_WRDATA_4(30),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_93);
  x_grlfpc2_0_wrdata_0_0_27x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(27),
    I1 => GRLFPC2_0_COMB_WRDATA_4(27),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_90);
  x_grlfpc2_0_wrdata_0_0_1x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(1),
    I1 => GRLFPC2_0_COMB_WRDATA_4(1),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_64);
  x_grlfpc2_0_comb_rs1_1_2_am_0x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_d_inst(14),
    I1 => GRLFPC2_0_R_A_RS1(0),
    I2 => holdn,
    O => N_12274);
  x_grlfpc2_0_comb_rs1_1_2_bm_0x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => cpi_d_inst(25),
    I1 => GRLFPC2_0_RS1V_0_SQMUXA,
    O => N_12275);
  x_grlfpc2_0_comb_rs1_1_2_0x: MUXF5 port map (
      I0 => N_12274,
      I1 => N_12275,
      S => GRLFPC2_0_COMB_RS2_1_SN_N_2,
      O => GRLFPC2_0_COMB_RS1_1(0));
  x_grlfpc2_0_comb_rs1_1_0_am_4x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_d_inst(18),
    I1 => GRLFPC2_0_R_A_RS1(4),
    I2 => holdn,
    O => N_12276);
  x_grlfpc2_0_comb_rs1_1_0_bm_4x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => cpi_d_inst(29),
    I1 => GRLFPC2_0_RS1V_0_SQMUXA,
    O => N_12277);
  x_grlfpc2_0_comb_rs1_1_0_4x: MUXF5 port map (
      I0 => N_12276,
      I1 => N_12277,
      S => GRLFPC2_0_COMB_RS2_1_SN_N_2,
      O => GRLFPC2_0_COMB_RS1_1(4));
  x_grlfpc2_0_comb_rs1_1_0_am_3x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_d_inst(17),
    I1 => GRLFPC2_0_R_A_RS1(3),
    I2 => holdn,
    O => N_12278);
  x_grlfpc2_0_comb_rs1_1_0_bm_3x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => cpi_d_inst(28),
    I1 => GRLFPC2_0_RS1V_0_SQMUXA,
    O => N_12279);
  x_grlfpc2_0_comb_rs1_1_0_3x: MUXF5 port map (
      I0 => N_12278,
      I1 => N_12279,
      S => GRLFPC2_0_COMB_RS2_1_SN_N_2,
      O => GRLFPC2_0_COMB_RS1_1(3));
  x_grlfpc2_0_comb_rs1_1_0_am_2x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_d_inst(16),
    I1 => GRLFPC2_0_R_A_RS1(2),
    I2 => holdn,
    O => N_12280);
  x_grlfpc2_0_comb_rs1_1_0_bm_2x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => cpi_d_inst(27),
    I1 => GRLFPC2_0_RS1V_0_SQMUXA,
    O => N_12281);
  x_grlfpc2_0_comb_rs1_1_0_2x: MUXF5 port map (
      I0 => N_12280,
      I1 => N_12281,
      S => GRLFPC2_0_COMB_RS2_1_SN_N_2,
      O => GRLFPC2_0_COMB_RS1_1(2));
  x_grlfpc2_0_comb_rs1_1_2_am_1x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_d_inst(15),
    I1 => GRLFPC2_0_R_A_RS1(1),
    I2 => holdn,
    O => N_12282);
  x_grlfpc2_0_comb_rs1_1_2_bm_1x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => cpi_d_inst(26),
    I1 => GRLFPC2_0_RS1V_0_SQMUXA,
    O => N_12283);
  x_grlfpc2_0_comb_rs1_1_2_1x: MUXF5 port map (
      I0 => N_12282,
      I1 => N_12283,
      S => GRLFPC2_0_COMB_RS2_1_SN_N_2,
      O => GRLFPC2_0_COMB_RS1_1(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_86x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(27),
    I1 => GRLFPC2_0_FPO_FRAC(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_592);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_95x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(18),
    I1 => GRLFPC2_0_FPO_FRAC(20),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_583);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_81x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(32),
    I1 => GRLFPC2_0_FPO_FRAC(34),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_597);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_98x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(15),
    I1 => GRLFPC2_0_FPO_FRAC(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_580);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_106x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(7),
    I1 => GRLFPC2_0_FPO_FRAC(9),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_572);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_87x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(26),
    I1 => GRLFPC2_0_FPO_FRAC(28),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_591);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_85x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(28),
    I1 => GRLFPC2_0_FPO_FRAC(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_593);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_84x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(29),
    I1 => GRLFPC2_0_FPO_FRAC(31),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_594);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_96x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(17),
    I1 => GRLFPC2_0_FPO_FRAC(19),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_582);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_0x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_16x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(17),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_15x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(15),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(16),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_4x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(5),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_78x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(35),
    I1 => GRLFPC2_0_FPO_FRAC(37),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_600);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_45x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(45),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(46),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_am_44x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(44),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(46),
    O => N_12284);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_bm_44x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(45),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(47),
    O => N_12285);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_44x: MUXF5 port map (
      I0 => N_12284,
      I1 => N_12285,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_65x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(48),
    I1 => GRLFPC2_0_FPO_FRAC(50),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_613);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_61x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(52),
    I1 => GRLFPC2_0_FPO_FRAC(54),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_617);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_60x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(53),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_278,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_618);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_am_54x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(54),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(56),
    O => N_12286);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_bm_54x: LUT3 
  generic map(
    INIT => X"74"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(57),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(55),
    O => N_12287);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_54x: MUXF5 port map (
      I0 => N_12286,
      I1 => N_12287,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_47x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(47),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(48),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_0_46x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(46),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(47),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_83x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(30),
    I1 => GRLFPC2_0_FPO_FRAC(32),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_595);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_91x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(22),
    I1 => GRLFPC2_0_FPO_FRAC(24),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_587);
  x_grlfpc2_0_wrdata_0_0_52x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(20),
    I1 => GRLFPC2_0_COMB_WRDATA_4(52),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_115);
  x_grlfpc2_0_wrdata_0_0_49x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(17),
    I1 => GRLFPC2_0_COMB_WRDATA_4(49),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_112);
  x_grlfpc2_0_wrdata_0_0_48x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(16),
    I1 => GRLFPC2_0_COMB_WRDATA_4(48),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_111);
  x_grlfpc2_0_wrdata_0_0_45x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(13),
    I1 => GRLFPC2_0_COMB_WRDATA_4(45),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_108);
  x_grlfpc2_0_wrdata_0_0_35x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(3),
    I1 => GRLFPC2_0_COMB_WRDATA_4(35),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_98);
  x_grlfpc2_0_wrdata_0_0_20x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(20),
    I1 => GRLFPC2_0_COMB_WRDATA_4(20),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_83);
  x_grlfpc2_0_wrdata_0_0_17x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(17),
    I1 => GRLFPC2_0_COMB_WRDATA_4(17),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_80);
  x_grlfpc2_0_wrdata_0_0_16x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(16),
    I1 => GRLFPC2_0_COMB_WRDATA_4(16),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_79);
  x_grlfpc2_0_wrdata_0_0_13x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(13),
    I1 => GRLFPC2_0_COMB_WRDATA_4(13),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_76);
  x_grlfpc2_0_wrdata_0_0_3x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_lddata(3),
    I1 => GRLFPC2_0_COMB_WRDATA_4(3),
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA_1,
    O => GRLFPC2_0_N_66);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_55_CA_2_55x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(57),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(316),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1932);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_CA_3_54x: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(57),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(316),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1933);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notstickyinforsr_2_1: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1870,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_49_1_2_258x: LUT3 
  generic map(
    INIT => X"96"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_49_1_0(258),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_49_1_2(258));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_waitmulxff_notsampledwait_i: LUT4 
  generic map(
    INIT => X"37F7"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN17_WQSTSETS,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_56_1: LUT3 
  generic map(
    INIT => X"95"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1533,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(59),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_56_I_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_57_1: LUT4 
  generic map(
    INIT => X"56FC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(58),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(174),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_1(0),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_57_I_1);
  x_grlfpc2_0_comb_v_state_7_1x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_R_STATE(1),
    I1 => GRLFPC2_0_V_STATE_2_SQMUXA,
    O => GRLFPC2_0_COMB_V_STATE_7(1));
  x_grlfpc2_0_comb_rs1v_1_i: LUT4 
  generic map(
    INIT => X"04CC"
  )
  port map (
    I0 => cpi_d_inst(30),
    I1 => cpi_d_inst(31),
    I2 => GRLFPC2_0_N_764,
    I3 => GRLFPC2_0_UN1_WREN210_4_0,
    O => GRLFPC2_0_COMB_RS1V_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_startshft_un3_notresetorunimp: LUT3 
  generic map(
    INIT => X"54"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTDECODEDUNIMP,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(65),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(66),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTRESETORUNIMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_c_pxs_multiplexormulxff_result_0_0_5x: LUT3 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => N_2461,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(55),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT0(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_c_pxs_multiplexormulxff_result_0_0_6x: LUT3 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => N_2462,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(54),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT0(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_c_pxs_multiplexormulxff_result_0_0_7x: LUT3 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => N_2463,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(53),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT0(7));
  x_grlfpc2_0_I_185_0_am: LUT4 
  generic map(
    INIT => X"3200"
  )
  port map (
    I0 => cpi_d_inst(14),
    I1 => GRLFPC2_0_COMB_FPDECODE_MOV5,
    I2 => GRLFPC2_0_COMB_RSDECODE_RS1V2_0,
    I3 => GRLFPC2_0_MOV_7_SQMUXA_3,
    O => N_12288);
  x_grlfpc2_0_I_185_0_bm: LUT3 
  generic map(
    INIT => X"20"
  )
  port map (
    I0 => cpi_d_inst(14),
    I1 => GRLFPC2_0_COMB_FPDECODE_RS2D5,
    I2 => GRLFPC2_0_MOV_7_SQMUXA_3,
    O => N_12289);
  x_grlfpc2_0_I_185_0: MUXF5 port map (
      I0 => N_12288,
      I1 => N_12289,
      S => cpi_d_inst(19),
      O => GRLFPC2_0_N_631);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlcregxz_un17_inforcregsn: LUT4_L 
  generic map(
    INIT => X"9000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2276,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2281_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_UN17_INFORCREGSN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_startshft_un2_notdecodedunimp: LUT3 
  generic map(
    INIT => X"10"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTDECODEDUNIMP,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(64),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(66),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN2_NOTDECODEDUNIMP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_7: LUT4 
  generic map(
    INIT => X"59A6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(7),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_1(49),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_7_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_11: LUT4 
  generic map(
    INIT => X"59A6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(11),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(11),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_1(45),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_11_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_15: LUT4 
  generic map(
    INIT => X"59A6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(15),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(15),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_1(41),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_15_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_17: LUT4 
  generic map(
    INIT => X"59A6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(17),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_1(39),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_17_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_2: LUT4 
  generic map(
    INIT => X"59A6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_1(54),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_2_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_21: LUT4 
  generic map(
    INIT => X"59A6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(21),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_1(35),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_21_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_25: LUT4 
  generic map(
    INIT => X"59A6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(25),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(25),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_1(31),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_25_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_26: LUT4 
  generic map(
    INIT => X"59A6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(26),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(26),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_1(30),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_26_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_27: LUT4 
  generic map(
    INIT => X"59A6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(27),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(27),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_1(29),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_27_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_32: LUT4_L 
  generic map(
    INIT => X"956A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1557,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_32_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_3: LUT4 
  generic map(
    INIT => X"59A6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_1(53),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_3_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_36: LUT4 
  generic map(
    INIT => X"956A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1553,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(79),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_36_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_37: LUT4 
  generic map(
    INIT => X"956A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1552,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(78),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_37_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_38: LUT4 
  generic map(
    INIT => X"956A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1551,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(77),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_38_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_39: LUT4 
  generic map(
    INIT => X"956A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1550,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_39_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_40: LUT4_L 
  generic map(
    INIT => X"956A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1549,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_40_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_41: LUT4_L 
  generic map(
    INIT => X"956A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1548,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(74),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_41_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_43: LUT4 
  generic map(
    INIT => X"956A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1546,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(72),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_43_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_45: LUT4_L 
  generic map(
    INIT => X"956A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1544,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(70),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_45_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_46: LUT4 
  generic map(
    INIT => X"956A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1543,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(69),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_46_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_47: LUT4 
  generic map(
    INIT => X"956A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1542,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(68),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_47_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_50: LUT4 
  generic map(
    INIT => X"956A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1539,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(65),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_50_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_52: LUT4_L 
  generic map(
    INIT => X"956A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1537,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(63),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_52_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_33: LUT4_L 
  generic map(
    INIT => X"956A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1556,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(82),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_33_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_34: LUT4 
  generic map(
    INIT => X"956A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1555,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(81),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_34_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_35: LUT4_L 
  generic map(
    INIT => X"956A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1554,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(80),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_35_I);
  x_grlfpc2_0_comb_fpdecode_st_0: LUT4 
  generic map(
    INIT => X"0C8C"
  )
  port map (
    I0 => cpi_d_inst(21),
    I1 => GRLFPC2_0_COMB_FPDECODE_AFQ13,
    I2 => GRLFPC2_0_UN1_AFQ3_I,
    I3 => GRLFPC2_0_UN1_AFQ6_I,
    O => GRLFPC2_0_COMB_FPDECODE_ST);
  x_grlfpc2_0_un1_mov_1_sqmuxa: LUT4 
  generic map(
    INIT => X"002F"
  )
  port map (
    I0 => GRLFPC2_0_N_766,
    I1 => GRLFPC2_0_COMB_FPDECODE_MOV5,
    I2 => GRLFPC2_0_COMB_FPDECODE_MOV11,
    I3 => GRLFPC2_0_MOV_2_SQMUXA,
    O => GRLFPC2_0_N_757);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_5: LUT4 
  generic map(
    INIT => X"59A6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(5),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_1(51),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_5_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_54: LUT4 
  generic map(
    INIT => X"956A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1535,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(61),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_54_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_53: LUT4 
  generic map(
    INIT => X"59A6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(53),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(3),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_53_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_51: LUT4_L 
  generic map(
    INIT => X"956A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1538,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_51_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_49: LUT4_L 
  generic map(
    INIT => X"956A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1540,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_49_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un22_xzxbus_48: LUT4_L 
  generic map(
    INIT => X"956A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1541,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(67),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_48_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_checkovanddenorm_un20_notpossibleov_4: LUT4 
  generic map(
    INIT => X"8000"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(47),
    I1 => GRLFPC2_0_FPO_FRAC(48),
    I2 => GRLFPC2_0_FPO_FRAC(49),
    I3 => GRLFPC2_0_FPO_FRAC(50),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CHECKOVANDDENORM_UN20_NOTPOSSIBLEOV_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_checkovanddenorm_un20_notpossibleov_5: LUT4 
  generic map(
    INIT => X"8000"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(51),
    I1 => GRLFPC2_0_FPO_FRAC(52),
    I2 => GRLFPC2_0_FPO_FRAC(53),
    I3 => GRLFPC2_0_FPO_FRAC(54),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CHECKOVANDDENORM_UN20_NOTPOSSIBLEOV_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_28_0_0: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CONDMUXMULXFF_UN4_NOTSQRTLFTCC,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14(77),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_50_trfwwbasiccell_un443_ca_i: LUT2 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1936,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_7(50),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_UN443_CA_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un22_gen: LUT4 
  generic map(
    INIT => X"E000"
  )
  port map (
    I0 => N_8928,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_57_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SALSBS(0),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_1(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN22_GEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un30_gen: LUT4 
  generic map(
    INIT => X"C888"
  )
  port map (
    I0 => N_8928,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_57_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(3),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN30_GEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_47_trfwwbasiccell_un462_ca_i: LUT3 
  generic map(
    INIT => X"40"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1939,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_TEMP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_UN462_CA_I);
  x_grlfpc2_0_comb_un6_rs1v: LUT2 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RS1_1(0),
    I1 => GRLFPC2_0_COMB_RS1D_1,
    O => GRLFPC2_0_N_752);
  x_grlfpc2_0_comb_un1_rs1v: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RS1_1(0),
    I1 => GRLFPC2_0_COMB_RS1D_1,
    O => GRLFPC2_0_N_751);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_1_3_209: LUT4 
  generic map(
    INIT => X"2242"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(57),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(316),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => N_2362);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_temp_2_1_1x: LUT3 
  generic map(
    INIT => X"54"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1987,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SBLSBS_0(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_CIN,
    O => N_8929);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_tz_375x: LUT4 
  generic map(
    INIT => X"02C2"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(52),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELINITREMBIT,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(61),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_TZ(375));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_57: LUT4 
  generic map(
    INIT => X"3666"
  )
  port map (
    I0 => N_8928,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_57_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(3),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN22_NOTPROP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_selectdivmult_un86_divmultv_0: LUT4 
  generic map(
    INIT => X"010D"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(52),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELINITREMBIT,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(61),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_TZ(375));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_94_1: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_94_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1942,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_129_1(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_96_1: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_96_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1943,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_130_1(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_98_1: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_98_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1962,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_149_1(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_61_1: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_61_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1948,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_135_1(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_62_1: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_62_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1963,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_150_1(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_66_1: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_66_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1964,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_151_1(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_74_1: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_74_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1953,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_140_1(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_78_1: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_78_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1950,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_137_1(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_101_12x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1972,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_43(14),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_101(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_95_18x: LUT4 
  generic map(
    INIT => X"69A5"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1966,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_37(20),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_TEMP2_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_95(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_111_2x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1982,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_53(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_111(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_109_4x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1980,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_51(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_109(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_108_5x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1979,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_50(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_108(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_94_19x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1965,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_36(21),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_94(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_87_26x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1958,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_29(28),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_87(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_si_113_0x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1984,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_113_0(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_113(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_64_49x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1935,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_6(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_64(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_83_30x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1954,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_25(32),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_83(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_81_32x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1952,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_23(34),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_81(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_80_33x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1951,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_22(35),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_80(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_73_40x: LUT4 
  generic map(
    INIT => X"69A5"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1944,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_15(42),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_TEMP2_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_73(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_74_39x: LUT4 
  generic map(
    INIT => X"69A5"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1945,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_16(41),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_TEMP2_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_74(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_85_28x: LUT4 
  generic map(
    INIT => X"69A5"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1956,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_27(30),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_TEMP2_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_85(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_86_27x: LUT4 
  generic map(
    INIT => X"69A5"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1957,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_28(29),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_TEMP2_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_86(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_90_23x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1961,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_32(25),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_90(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_106_7x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1977,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_48(9),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_106(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_84_29x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1955,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_26(31),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_84(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_69_44x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1940,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_11(46),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_69(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_98_15x: LUT4 
  generic map(
    INIT => X"69A5"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1969,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_40(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_TEMP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_98(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_70_43x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1941,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_12(45),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_70(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_64_1: LUT4 
  generic map(
    INIT => X"6999"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_64_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1939,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_TEMP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_68(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_67_46x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1938,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_9(48),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_67(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_105_8x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1976,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_47(10),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_105(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_107_6x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1978,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_49(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_107(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_103_10x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1974,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_45(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_103(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_SBLSBs_0x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1987,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SBLSBS_0(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SBLSBS(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_SBLSBs_1_1x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1985,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SBLSBS_1_0(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SBLSBS_1(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_100_13x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1971,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_42(15),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_100(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_102_11x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1973,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_44(13),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_102(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_99_14x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1970,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_41(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_99(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_97_16x: LUT4 
  generic map(
    INIT => X"69A5"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1968,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_39(18),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_18_TRFWWBASICCELL_TEMP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_97(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_104_9x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1975,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_46(11),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_104(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_104_1: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_104_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1981,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_168_1(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_100_1: LUT4 
  generic map(
    INIT => X"6999"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_100_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1967,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_19_TRFWWBASICCELL_TEMP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_154_1(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_75_38x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1946,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_17(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_75(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_76_37x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1947,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_18(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_76(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_78_35x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1949,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_20(37),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_78(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_89_24x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1960,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_31(26),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_89(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_88_1: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_88_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1959,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_88(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_65_48x: LUT4 
  generic map(
    INIT => X"69A5"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1936,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_7(50),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_TEMP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_65(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_66_47x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1937,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_8(49),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_66(47));
  x_grlfpc2_0_I_237_0: LUT4 
  generic map(
    INIT => X"9382"
  )
  port map (
    I0 => cpi_d_inst(19),
    I1 => cpi_d_inst(20),
    I2 => cpi_d_inst(30),
    I3 => GRLFPC2_0_N_674,
    O => GRLFPC2_0_I_237_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notstickyinforsr_2_2: LUT4_L 
  generic map(
    INIT => X"080A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_2_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN24_SHDVAR,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_UN57_SHDVAR,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(2),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_2_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_NE_7: LUT4 
  generic map(
    INIT => X"0100"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_7,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_8,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_9,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_NE_4,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_NE_7);
  x_grlfpc2_0_comb_v_state_7_iv_0x: LUT4 
  generic map(
    INIT => X"8CAF"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_I_V6,
    I1 => GRLFPC2_0_R_STATE(0),
    I2 => GRLFPC2_0_V_STATE_1_SQMUXA_3_0,
    I3 => GRLFPC2_0_V_STATE_2_SQMUXA,
    O => GRLFPC2_0_COMB_V_STATE_7(0));
  x_grlfpc2_0_I_196: LUT2 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => cpi_d_inst(30),
    I1 => GRLFPC2_0_N_631,
    O => GRLFPC2_0_N_636);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un2_notabortwb: LUT4 
  generic map(
    INIT => X"AAA8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14(77),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(77),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_se_0_4x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(4),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_se_0_6x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_se_0_10x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(10),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(11),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_se_0_11x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(11),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_se_0_16x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(16),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_se_0_18x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(18),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(19),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_se_0_20x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(20),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(21),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_se_0_21x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(22),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_se_0_22x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(22),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(23),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_se_0_23x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(24),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_se_0_24x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(24),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(25),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_se_0_26x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(26),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(27),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_se_0_27x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(27),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(28),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_se_0_28x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(28),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_se_0_30x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(31),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_se_0_31x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(31),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(32),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_se_0_33x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(33),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(34),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_se_0_36x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(36),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(37),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_se_0_46x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(46),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(47),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_pxs_multiplexormulxff_result_0_0_0_3x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => N_2459,
    I1 => cpi_d_inst(11),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_71,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_76);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_14_0_0_am: LUT4 
  generic map(
    INIT => X"C939"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(244),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(48),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(52),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(12),
    O => N_12290);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_14_0_0_bm: LUT4 
  generic map(
    INIT => X"5AC3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN42_CONDITIONAL,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_CONDITIONAL(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(48),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(52),
    O => N_12291);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_14_0_0: MUXF5 port map (
      I0 => N_12290,
      I1 => N_12291,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(51),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_360);
  x_grlfpc2_0_comb_v_i_res_1_0_am_29x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_FRAC(32),
    I2 => GRLFPC2_0_R_I_RES(29),
    O => N_12292);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_29x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(0),
    I2 => rfo2_data2(0),
    O => N_12293);
  x_grlfpc2_0_comb_v_i_res_1_0_29x: MUXF5 port map (
      I0 => N_12292,
      I1 => N_12293,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(29));
  x_grlfpc2_0_comb_v_i_res_1_0_am_30x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_FRAC(33),
    I2 => GRLFPC2_0_R_I_RES(30),
    O => N_12294);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_30x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(1),
    I2 => rfo2_data2(1),
    O => N_12295);
  x_grlfpc2_0_comb_v_i_res_1_0_30x: MUXF5 port map (
      I0 => N_12294,
      I1 => N_12295,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(30));
  x_grlfpc2_0_comb_v_i_res_1_0_am_31x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_FRAC(34),
    I2 => GRLFPC2_0_R_I_RES(31),
    O => N_12296);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_31x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(2),
    I2 => rfo2_data2(2),
    O => N_12297);
  x_grlfpc2_0_comb_v_i_res_1_0_31x: MUXF5 port map (
      I0 => N_12296,
      I1 => N_12297,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(31));
  x_grlfpc2_0_comb_v_i_res_1_0_am_34x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_FRAC(37),
    I2 => GRLFPC2_0_R_I_RES(34),
    O => N_12298);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_34x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(5),
    I2 => rfo2_data2(5),
    O => N_12299);
  x_grlfpc2_0_comb_v_i_res_1_0_34x: MUXF5 port map (
      I0 => N_12298,
      I1 => N_12299,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(34));
  x_grlfpc2_0_comb_v_i_res_1_0_am_36x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_FRAC(39),
    I2 => GRLFPC2_0_R_I_RES(36),
    O => N_12300);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_36x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(7),
    I2 => rfo2_data2(7),
    O => N_12301);
  x_grlfpc2_0_comb_v_i_res_1_0_36x: MUXF5 port map (
      I0 => N_12300,
      I1 => N_12301,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(36));
  x_grlfpc2_0_comb_v_i_res_1_0_am_37x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_FRAC(40),
    I2 => GRLFPC2_0_R_I_RES(37),
    O => N_12302);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_37x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(8),
    I2 => rfo2_data2(8),
    O => N_12303);
  x_grlfpc2_0_comb_v_i_res_1_0_37x: MUXF5 port map (
      I0 => N_12302,
      I1 => N_12303,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(37));
  x_grlfpc2_0_comb_v_i_res_1_0_am_38x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_FRAC(41),
    I2 => GRLFPC2_0_R_I_RES(38),
    O => N_12304);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_38x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(9),
    I2 => rfo2_data2(9),
    O => N_12305);
  x_grlfpc2_0_comb_v_i_res_1_0_38x: MUXF5 port map (
      I0 => N_12304,
      I1 => N_12305,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(38));
  x_grlfpc2_0_comb_v_i_res_1_0_am_39x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_FRAC(42),
    I2 => GRLFPC2_0_R_I_RES(39),
    O => N_12306);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_39x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(10),
    I2 => rfo2_data2(10),
    O => N_12307);
  x_grlfpc2_0_comb_v_i_res_1_0_39x: MUXF5 port map (
      I0 => N_12306,
      I1 => N_12307,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(39));
  x_grlfpc2_0_comb_v_i_res_1_0_am_40x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_FRAC(43),
    I2 => GRLFPC2_0_R_I_RES(40),
    O => N_12308);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_40x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(11),
    I2 => rfo2_data2(11),
    O => N_12309);
  x_grlfpc2_0_comb_v_i_res_1_0_40x: MUXF5 port map (
      I0 => N_12308,
      I1 => N_12309,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(40));
  x_grlfpc2_0_comb_v_i_res_1_0_am_41x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_FRAC(44),
    I2 => GRLFPC2_0_R_I_RES(41),
    O => N_12310);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_41x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(12),
    I2 => rfo2_data2(12),
    O => N_12311);
  x_grlfpc2_0_comb_v_i_res_1_0_41x: MUXF5 port map (
      I0 => N_12310,
      I1 => N_12311,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(41));
  x_grlfpc2_0_comb_v_i_res_1_0_am_42x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_FRAC(45),
    I2 => GRLFPC2_0_R_I_RES(42),
    O => N_12312);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_42x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(13),
    I2 => rfo2_data2(13),
    O => N_12313);
  x_grlfpc2_0_comb_v_i_res_1_0_42x: MUXF5 port map (
      I0 => N_12312,
      I1 => N_12313,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(42));
  x_grlfpc2_0_comb_v_i_res_1_0_am_43x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_FRAC(46),
    I2 => GRLFPC2_0_R_I_RES(43),
    O => N_12314);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_43x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(14),
    I2 => rfo2_data2(14),
    O => N_12315);
  x_grlfpc2_0_comb_v_i_res_1_0_43x: MUXF5 port map (
      I0 => N_12314,
      I1 => N_12315,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(43));
  x_grlfpc2_0_comb_v_i_res_1_0_am_44x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_FRAC(47),
    I2 => GRLFPC2_0_R_I_RES(44),
    O => N_12316);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_44x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(15),
    I2 => rfo2_data2(15),
    O => N_12317);
  x_grlfpc2_0_comb_v_i_res_1_0_44x: MUXF5 port map (
      I0 => N_12316,
      I1 => N_12317,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(44));
  x_grlfpc2_0_comb_v_i_res_1_0_am_45x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_FRAC(48),
    I2 => GRLFPC2_0_R_I_RES(45),
    O => N_12318);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_45x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(16),
    I2 => rfo2_data2(16),
    O => N_12319);
  x_grlfpc2_0_comb_v_i_res_1_0_45x: MUXF5 port map (
      I0 => N_12318,
      I1 => N_12319,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(45));
  x_grlfpc2_0_comb_v_i_res_1_0_am_46x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_FRAC(49),
    I2 => GRLFPC2_0_R_I_RES(46),
    O => N_12320);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_46x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(17),
    I2 => rfo2_data2(17),
    O => N_12321);
  x_grlfpc2_0_comb_v_i_res_1_0_46x: MUXF5 port map (
      I0 => N_12320,
      I1 => N_12321,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(46));
  x_grlfpc2_0_comb_v_i_res_1_0_am_47x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_FRAC(50),
    I2 => GRLFPC2_0_R_I_RES(47),
    O => N_12322);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_47x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(18),
    I2 => rfo2_data2(18),
    O => N_12323);
  x_grlfpc2_0_comb_v_i_res_1_0_47x: MUXF5 port map (
      I0 => N_12322,
      I1 => N_12323,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(47));
  x_grlfpc2_0_comb_v_i_res_1_0_am_49x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_FRAC(52),
    I2 => GRLFPC2_0_R_I_RES(49),
    O => N_12324);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_49x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(20),
    I2 => rfo2_data2(20),
    O => N_12325);
  x_grlfpc2_0_comb_v_i_res_1_0_49x: MUXF5 port map (
      I0 => N_12324,
      I1 => N_12325,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(49));
  x_grlfpc2_0_comb_v_i_res_1_0_am_50x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_FRAC(53),
    I2 => GRLFPC2_0_R_I_RES(50),
    O => N_12326);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_50x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(21),
    I2 => rfo2_data2(21),
    O => N_12327);
  x_grlfpc2_0_comb_v_i_res_1_0_50x: MUXF5 port map (
      I0 => N_12326,
      I1 => N_12327,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(50));
  x_grlfpc2_0_comb_v_i_res_1_0_am_51x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_FRAC(54),
    I2 => GRLFPC2_0_R_I_RES(51),
    O => N_12328);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_51x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(22),
    I2 => rfo2_data2(22),
    O => N_12329);
  x_grlfpc2_0_comb_v_i_res_1_0_51x: MUXF5 port map (
      I0 => N_12328,
      I1 => N_12329,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(51));
  x_grlfpc2_0_wrdata_0_0x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(0),
    I1 => GRLFPC2_0_N_63,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(0));
  x_grlfpc2_0_wrdata_1_1x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(1),
    I1 => GRLFPC2_0_N_64,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(1));
  x_grlfpc2_0_wrdata_0_2x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(2),
    I1 => GRLFPC2_0_N_65,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(2));
  x_grlfpc2_0_wrdata_1_3x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(3),
    I1 => GRLFPC2_0_N_66,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(3));
  x_grlfpc2_0_wrdata_0_4x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(4),
    I1 => GRLFPC2_0_N_67,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(4));
  x_grlfpc2_0_wrdata_0_5x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(5),
    I1 => GRLFPC2_0_N_68,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(5));
  x_grlfpc2_0_wrdata_0_6x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(6),
    I1 => GRLFPC2_0_N_69,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(6));
  x_grlfpc2_0_wrdata_0_7x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(7),
    I1 => GRLFPC2_0_N_70,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(7));
  x_grlfpc2_0_wrdata_0_8x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(8),
    I1 => GRLFPC2_0_N_71,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(8));
  x_grlfpc2_0_wrdata_0_9x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(9),
    I1 => GRLFPC2_0_N_72,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(9));
  x_grlfpc2_0_wrdata_0_10x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(10),
    I1 => GRLFPC2_0_N_73,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(10));
  x_grlfpc2_0_wrdata_0_11x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(11),
    I1 => GRLFPC2_0_N_74,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(11));
  x_grlfpc2_0_wrdata_0_12x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(12),
    I1 => GRLFPC2_0_N_75,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(12));
  x_grlfpc2_0_wrdata_0_14x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(14),
    I1 => GRLFPC2_0_N_77,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(14));
  x_grlfpc2_0_wrdata_0_15x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(15),
    I1 => GRLFPC2_0_N_78,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(15));
  x_grlfpc2_0_wrdata_0_18x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(18),
    I1 => GRLFPC2_0_N_81,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(18));
  x_grlfpc2_0_wrdata_0_19x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(19),
    I1 => GRLFPC2_0_N_82,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(19));
  x_grlfpc2_0_wrdata_0_21x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(21),
    I1 => GRLFPC2_0_N_84,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(21));
  x_grlfpc2_0_wrdata_0_22x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(22),
    I1 => GRLFPC2_0_N_85,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(22));
  x_grlfpc2_0_wrdata_0_23x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(23),
    I1 => GRLFPC2_0_N_86,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(23));
  x_grlfpc2_0_wrdata_0_24x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(24),
    I1 => GRLFPC2_0_N_87,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(24));
  x_grlfpc2_0_wrdata_0_25x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(25),
    I1 => GRLFPC2_0_N_88,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(25));
  x_grlfpc2_0_wrdata_0_26x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(26),
    I1 => GRLFPC2_0_N_89,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(26));
  x_grlfpc2_0_wrdata_0_28x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(28),
    I1 => GRLFPC2_0_N_91,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(28));
  x_grlfpc2_0_wrdata_0_29x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(29),
    I1 => GRLFPC2_0_N_92,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(29));
  x_grlfpc2_0_wrdata_0_31x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(31),
    I1 => GRLFPC2_0_N_94,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(31));
  x_grlfpc2_0_wrdata_0_32x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(0),
    I1 => GRLFPC2_0_N_95,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(0));
  x_grlfpc2_0_wrdata_0_34x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(2),
    I1 => GRLFPC2_0_N_97,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(2));
  x_grlfpc2_0_wrdata_0_36x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(4),
    I1 => GRLFPC2_0_N_99,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(4));
  x_grlfpc2_0_wrdata_0_37x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(5),
    I1 => GRLFPC2_0_N_100,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(5));
  x_grlfpc2_0_wrdata_0_38x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(6),
    I1 => GRLFPC2_0_N_101,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(6));
  x_grlfpc2_0_wrdata_0_39x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(7),
    I1 => GRLFPC2_0_N_102,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(7));
  x_grlfpc2_0_wrdata_0_40x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(8),
    I1 => GRLFPC2_0_N_103,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(8));
  x_grlfpc2_0_wrdata_0_41x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(9),
    I1 => GRLFPC2_0_N_104,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(9));
  x_grlfpc2_0_wrdata_0_42x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(10),
    I1 => GRLFPC2_0_N_105,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(10));
  x_grlfpc2_0_wrdata_0_43x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(11),
    I1 => GRLFPC2_0_N_106,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(11));
  x_grlfpc2_0_wrdata_0_44x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(12),
    I1 => GRLFPC2_0_N_107,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(12));
  x_grlfpc2_0_wrdata_0_46x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(14),
    I1 => GRLFPC2_0_N_109,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(14));
  x_grlfpc2_0_wrdata_0_47x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(15),
    I1 => GRLFPC2_0_N_110,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(15));
  x_grlfpc2_0_wrdata_0_50x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(18),
    I1 => GRLFPC2_0_N_113,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(18));
  x_grlfpc2_0_wrdata_0_51x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(19),
    I1 => GRLFPC2_0_N_114,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(19));
  x_grlfpc2_0_wrdata_0_53x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(21),
    I1 => GRLFPC2_0_N_116,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(21));
  x_grlfpc2_0_wrdata_0_54x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(22),
    I1 => GRLFPC2_0_N_117,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(22));
  x_grlfpc2_0_wrdata_0_55x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(23),
    I1 => GRLFPC2_0_N_118,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(23));
  x_grlfpc2_0_wrdata_0_56x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(24),
    I1 => GRLFPC2_0_N_119,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(24));
  x_grlfpc2_0_wrdata_0_57x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(25),
    I1 => GRLFPC2_0_N_120,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(25));
  x_grlfpc2_0_wrdata_0_58x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(26),
    I1 => GRLFPC2_0_N_121,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(26));
  x_grlfpc2_0_wrdata_0_60x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(28),
    I1 => GRLFPC2_0_N_123,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(28));
  x_grlfpc2_0_wrdata_0_61x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(29),
    I1 => GRLFPC2_0_N_124,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(29));
  x_grlfpc2_0_wrdata_1_62x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(30),
    I1 => GRLFPC2_0_N_125,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(30));
  x_grlfpc2_0_wrdata_1_59x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(27),
    I1 => GRLFPC2_0_N_122,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(27));
  x_grlfpc2_0_wrdata_1_33x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(1),
    I1 => GRLFPC2_0_N_96,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(1));
  x_grlfpc2_0_wrdata_1_30x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(30),
    I1 => GRLFPC2_0_N_93,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(30));
  x_grlfpc2_0_wrdata_1_27x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(27),
    I1 => GRLFPC2_0_N_90,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_c_pxs_multiplexormulxff_result_0_0_0x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => N_2456,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT0(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_se_0_17x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(17),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(18),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_se_0_25x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(25),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(26),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_se_0_37x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(37),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(38),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(37));
  x_grlfpc2_0_comb_v_i_res_1_0_am_48x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => GRLFPC2_0_FPO_FRAC(51),
    I2 => GRLFPC2_0_R_I_RES(48),
    O => N_12330);
  x_grlfpc2_0_comb_v_i_res_1_0_bm_48x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_N_771,
    I1 => rfo1_data2(19),
    I2 => rfo2_data2(19),
    O => N_12331);
  x_grlfpc2_0_comb_v_i_res_1_0_48x: MUXF5 port map (
      I0 => N_12330,
      I1 => N_12331,
      S => GRLFPC2_0_COMB_UN2_HOLDN,
      O => GRLFPC2_0_COMB_V_I_RES_1(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_se_0_2x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_se_0_1x: LUT3 
  generic map(
    INIT => X"35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(1));
  x_grlfpc2_0_rs1_1_0_1x: LUT3 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => cpi_dbg_addr(1),
    I1 => cpi_dbg_enable,
    I2 => GRLFPC2_0_COMB_RS1_1(1),
    O => RFI2_RD1ADDR_0_INT_5_INT_17);
  x_grlfpc2_0_rs1_1_0_2x: LUT3 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => cpi_dbg_addr(2),
    I1 => cpi_dbg_enable,
    I2 => GRLFPC2_0_COMB_RS1_1(2),
    O => RFI2_RD1ADDR_1_INT_6_INT_18);
  x_grlfpc2_0_rs1_1_0_3x: LUT3 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => cpi_dbg_addr(3),
    I1 => cpi_dbg_enable,
    I2 => GRLFPC2_0_COMB_RS1_1(3),
    O => RFI2_RD1ADDR_2_INT_7_INT_19);
  x_grlfpc2_0_rs1_1_0_4x: LUT3 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => cpi_dbg_addr(4),
    I1 => cpi_dbg_enable,
    I2 => GRLFPC2_0_COMB_RS1_1(4),
    O => RFI2_RD1ADDR_3_INT_8_INT_20);
  x_grlfpc2_0_wrdata_1_52x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(20),
    I1 => GRLFPC2_0_N_115,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(20));
  x_grlfpc2_0_wrdata_1_49x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(17),
    I1 => GRLFPC2_0_N_112,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(17));
  x_grlfpc2_0_wrdata_1_48x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(16),
    I1 => GRLFPC2_0_N_111,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(16));
  x_grlfpc2_0_wrdata_1_45x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(13),
    I1 => GRLFPC2_0_N_108,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(13));
  x_grlfpc2_0_wrdata_1_35x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(3),
    I1 => GRLFPC2_0_N_98,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi1_wrdata(3));
  x_grlfpc2_0_wrdata_1_20x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(20),
    I1 => GRLFPC2_0_N_83,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(20));
  x_grlfpc2_0_wrdata_1_17x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(17),
    I1 => GRLFPC2_0_N_80,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(17));
  x_grlfpc2_0_wrdata_1_16x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(16),
    I1 => GRLFPC2_0_N_79,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(16));
  x_grlfpc2_0_wrdata_1_13x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(13),
    I1 => GRLFPC2_0_N_76,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    O => rfi2_wrdata(13));
  x_grlfpc2_0_comb_v_fsr_cexc_1_iv_0_2x: LUT4 
  generic map(
    INIT => X"553F"
  )
  port map (
    I0 => cpi_dbg_data(2),
    I1 => GRLFPC2_0_COMB_MEXC_1(2),
    I2 => GRLFPC2_0_COMB_V_I_V6,
    I3 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
    O => GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_0(2));
  x_grlfpc2_0_comb_v_fsr_cexc_1_iv_0_0x: LUT4 
  generic map(
    INIT => X"553F"
  )
  port map (
    I0 => cpi_dbg_data(0),
    I1 => GRLFPC2_0_COMB_MEXC_1(0),
    I2 => GRLFPC2_0_COMB_V_I_V6,
    I3 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
    O => GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_0(0));
  x_grlfpc2_0_comb_v_fsr_cexc_1_iv_0_3x: LUT4 
  generic map(
    INIT => X"553F"
  )
  port map (
    I0 => cpi_dbg_data(3),
    I1 => GRLFPC2_0_COMB_MEXC_1(3),
    I2 => GRLFPC2_0_COMB_V_I_V6,
    I3 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
    O => GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_0(3));
  x_grlfpc2_0_comb_v_fsr_cexc_1_iv_0_1x: LUT4 
  generic map(
    INIT => X"553F"
  )
  port map (
    I0 => cpi_dbg_data(1),
    I1 => GRLFPC2_0_COMB_MEXC_1(1),
    I2 => GRLFPC2_0_COMB_V_I_V6,
    I3 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
    O => GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_0(1));
  x_grlfpc2_0_comb_v_fsr_cexc_1_iv_0_4x: LUT4 
  generic map(
    INIT => X"553F"
  )
  port map (
    I0 => cpi_dbg_data(4),
    I1 => GRLFPC2_0_COMB_MEXC_1(4),
    I2 => GRLFPC2_0_COMB_V_I_V6,
    I3 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
    O => GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_0(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_1: LUT4 
  generic map(
    INIT => X"0012"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN20_XZXBUS(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_3: LUT4_L 
  generic map(
    INIT => X"8448"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1559,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_35_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(30),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_6: LUT4 
  generic map(
    INIT => X"8448"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1575,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_3_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(14),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_11: LUT4_L 
  generic map(
    INIT => X"8448"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1577,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_15_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(12),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_11);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_13: LUT4 
  generic map(
    INIT => X"8448"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1585,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_17_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(4),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_13);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_14: LUT4 
  generic map(
    INIT => X"8448"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1571,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_49_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(18),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_14);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_15: LUT4 
  generic map(
    INIT => X"8448"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1569,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_27_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(20),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_15);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_16: LUT4 
  generic map(
    INIT => X"8448"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1534,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_33_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(55),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_16);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_17: LUT4_L 
  generic map(
    INIT => X"8448"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1560,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_51_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(29),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_17);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_19: LUT4_L 
  generic map(
    INIT => X"8448"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1567,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_48_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(22),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_19);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_21: LUT4 
  generic map(
    INIT => X"8448"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1580,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_11_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(9),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_21);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_22: LUT4 
  generic map(
    INIT => X"8448"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1583,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_45_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(6),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_22);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_23: LUT4 
  generic map(
    INIT => X"8448"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1576,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_32_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(13),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_23);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_24: LUT4 
  generic map(
    INIT => X"8448"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1565,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_21_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(24),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_24);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_25: LUT4_L 
  generic map(
    INIT => X"8448"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1561,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_41_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(28),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_25);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_27: LUT4_L 
  generic map(
    INIT => X"8448"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1581,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_40_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(8),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_27);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_29: LUT4 
  generic map(
    INIT => X"8448"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1579,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_52_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(10),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_29);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_62_51x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1933,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_62_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_62(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_temp_2_1x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1987,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SBLSBS_0(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_2_I(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_63_50x: LUT4 
  generic map(
    INIT => X"9669"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1934,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_CIN_2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_114_1_1_0(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_63(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_feedback_0_2x: LUT4 
  generic map(
    INIT => X"7340"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(54),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN18_FEEDBACK,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_0(9),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(58),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_47_CA_67_0_47x: LUT4 
  generic map(
    INIT => X"A222"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_64_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1939,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_TEMP2,
    O => N_8863);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_50_CA_64_0_50x: LUT4 
  generic map(
    INIT => X"C400"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1936,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_7(50),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_TEMP2,
    O => N_8825);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_selectdivmult_un86_divmultv: LUT3 
  generic map(
    INIT => X"20"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_TZ(375),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SELECTDIVMULT_UN86_DIVMULTV);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_si_58_1_56x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1932,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_114_1_1_0(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_58_1(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_divmultv_0_a2_0_0x: LUT4 
  generic map(
    INIT => X"4000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(2),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(3),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2298);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_62_0: LUT4_L 
  generic map(
    INIT => X"9669"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_62_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1963,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_CIN,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_CIN_1,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_62_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_120_1_49x: LUT4 
  generic map(
    INIT => X"9669"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1933,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_62_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_CIN_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_120_1(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlcregxz_xzcregloaden_0_0_a2: LUT2 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_pxs_multiplexormulxff_result_0_sn_m4_i: LUT3 
  generic map(
    INIT => X"0E"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14(77),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTRESETORUNIMP,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1646);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlaregexp_exparegloaden_1: LUT2 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_1(68),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLOADEN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_un4_togglesig: LUT2 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(20),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN4_TOGGLESIG);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xztregloaden: LUT2 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_rndmodeselect_un1_temp: LUT2 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(21),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN1_TEMP);
  x_grlfpc2_0_comb_ccwr4_1: LUT4 
  generic map(
    INIT => X"0200"
  )
  port map (
    I0 => GRLFPC2_0_N_789,
    I1 => GRLFPC2_0_COMB_V_STATE_7(0),
    I2 => GRLFPC2_0_COMB_V_STATE_7(1),
    I3 => GRLFPC2_0_R_I_V,
    O => GRLFPC2_0_COMB_CCWR4_1);
  x_grlfpc2_0_comb_lockgen_locki_sn_m1_e: LUT4 
  generic map(
    INIT => X"1011"
  )
  port map (
    I0 => cpi_d_cnt(0),
    I1 => cpi_d_cnt(1),
    I2 => GRLFPC2_0_COMB_FPDECODE_ST,
    I3 => GRLFPC2_0_COMB_SEQERR_UN7_OP_I,
    O => GRLFPC2_0_COMB_LOCKGEN_LOCKI_SN_N_10);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_31: LUT4 
  generic map(
    INIT => X"9000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1573,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_16_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_26_I,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_27,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_31);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_32: LUT4 
  generic map(
    INIT => X"9000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1545,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_44_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_50_I,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_25,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_32);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_36: LUT4 
  generic map(
    INIT => X"9000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1570,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_19_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_25_I,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_17,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_36);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_39: LUT4 
  generic map(
    INIT => X"8400"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1566,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_2_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_23_0,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_11,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_39);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_40: LUT4 
  generic map(
    INIT => X"8000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_7_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_38_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_46_I,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_54_I,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_40);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_41: LUT4_L 
  generic map(
    INIT => X"8000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_34_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_36_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_47_I,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_53_I,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_41);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_43: LUT4 
  generic map(
    INIT => X"8400"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1547,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_37_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_42_0,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_43);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_un2_notabortwb_i: LUT4 
  generic map(
    INIT => X"5557"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14(77),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(77),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_notsrres_m_0_29x: LUT4 
  generic map(
    INIT => X"5044"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(30),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_notsrres_m_0_7x: LUT4 
  generic map(
    INIT => X"5044"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(8),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_notsrres_m_0_39x: LUT4 
  generic map(
    INIT => X"5044"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(40),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_notsrres_m_0_19x: LUT4 
  generic map(
    INIT => X"5044"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(19),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(20),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_notsrres_m_0_15x: LUT4 
  generic map(
    INIT => X"5044"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(15),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(16),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_notsrres_m_0_13x: LUT4 
  generic map(
    INIT => X"5044"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(13),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(14),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_notsrres_m_0_9x: LUT4 
  generic map(
    INIT => X"5044"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(9),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(10),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_notsrres_m_0_8x: LUT4 
  generic map(
    INIT => X"5044"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(9),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_notsrres_m_0_35x: LUT4 
  generic map(
    INIT => X"5044"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(35),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(36),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_notsrres_m_0_34x: LUT4 
  generic map(
    INIT => X"5044"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(34),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(35),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_notsrres_m_0_3x: LUT4 
  generic map(
    INIT => X"5044"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(4),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_notsrres_m_0_47x: LUT4 
  generic map(
    INIT => X"5044"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(47),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(48),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_notsrres_m_0_45x: LUT4 
  generic map(
    INIT => X"5044"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(45),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(46),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_notsrres_m_0_44x: LUT4 
  generic map(
    INIT => X"5044"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(44),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(45),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_notsrres_m_0_43x: LUT4 
  generic map(
    INIT => X"5044"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(43),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(44),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_notsrres_m_0_42x: LUT4 
  generic map(
    INIT => X"5044"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(43),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_notsrres_m_0_41x: LUT4 
  generic map(
    INIT => X"5044"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(41),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(42),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_notsrres_m_0_40x: LUT4 
  generic map(
    INIT => X"5044"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(41),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_notsrres_m_0_5x: LUT4 
  generic map(
    INIT => X"5044"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(6),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_notsrres_m_0_38x: LUT4 
  generic map(
    INIT => X"5044"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(38),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(39),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_notsrres_m_0_32x: LUT4 
  generic map(
    INIT => X"5044"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(32),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(33),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_busymulxff_un2_temp_1_0: LUT4 
  generic map(
    INIT => X"1000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_14(77),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN2_NOTDECODEDUNIMP,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(68),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(70),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_BUSYMULXFF_UN2_TEMP_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_122: LUT4 
  generic map(
    INIT => X"2DB4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1987,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SBLSBS_0(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SBLSBS_1(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN35_NOTPROP);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_46_CA_68_46x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1940,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_11(46),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1880);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_53_CA_61_53x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1933,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_62_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1873);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_CA_60_54x: LUT4 
  generic map(
    INIT => X"B22B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1932,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_CIN_3,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_114_1_1_0(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1872);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_55_CA_59_55x: LUT4 
  generic map(
    INIT => X"B22B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1932,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_CIN_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_CIN_3,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_114_1_1_0(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1871);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_33_CA_81_33x: LUT3 
  generic map(
    INIT => X"4D"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_74_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1953,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1893);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_36_CA_78_36x: LUT3 
  generic map(
    INIT => X"4D"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_78_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1950,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1890);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_38_CA_76_38x: LUT3 
  generic map(
    INIT => X"4D"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_61_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1948,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1888);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_40_CA_74_40x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1946,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_17(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1886);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_42_CA_72_42x: LUT4 
  generic map(
    INIT => X"2BAF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1944,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_15(42),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_TEMP2_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1884);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_43_CA_71_43x: LUT3 
  generic map(
    INIT => X"4D"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_96_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1943,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1883);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_44_CA_70_44x: LUT3 
  generic map(
    INIT => X"4D"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_94_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1942,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1882);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_20_CA_94_20x: LUT4 
  generic map(
    INIT => X"2BAF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1966,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_37(20),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_TEMP2_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1906);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_22_CA_92_22x: LUT3 
  generic map(
    INIT => X"4D"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_66_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1964,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1904);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_CA_91_23x: LUT3 
  generic map(
    INIT => X"4D"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_62_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1963,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1903);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_CA_90_24x: LUT3 
  generic map(
    INIT => X"4D"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_98_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1962,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1902);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_29_CA_85_29x: LUT4 
  generic map(
    INIT => X"2BAF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1957,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_28(29),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_TEMP2_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1897);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_CA_111_3x: LUT3 
  generic map(
    INIT => X"4D"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_13_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1983,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1923);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_5_CA_109_5x: LUT3 
  generic map(
    INIT => X"4D"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_104_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1981,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1921);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_27_CA_87_27x: LUT3 
  generic map(
    INIT => X"4D"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_88_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1959,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1899);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_21_CA_93_21x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1965,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_36(21),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1905);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_CA_107_7x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1979,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_50(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1919);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_6_CA_108_6x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1980,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_51(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1920);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_CA_110_4x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1982,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_53(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1922);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_41_CA_73_41x: LUT4 
  generic map(
    INIT => X"2BAF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1945,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_16(41),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_TEMP2_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1885);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_35_CA_79_35x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1951,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_22(35),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1891);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_34_CA_80_34x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1952,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_23(34),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1892);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_31_CA_83_31x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1955,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_26(31),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1895);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_52_CA_62_52x: LUT4 
  generic map(
    INIT => X"B22B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1934,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_CIN_2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_114_1_1_0(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1874);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_51_CA_63_51x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1935,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_6(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1875);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_48_CA_66_48x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1938,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_9(48),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1878);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_CA_112_2x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1984,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_113_0(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1924);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_25_CA_89_25x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1961,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_32(25),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1901);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_28_CA_86_28x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1958,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_29(28),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1898);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_30_CA_84_30x: LUT4 
  generic map(
    INIT => X"2BAF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1956,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_27(30),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_TEMP2_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1896);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_CA_105_9x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1977,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_48(9),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1917);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_12_CA_102_12x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1974,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_45(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1914);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_CA_103_11x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1975,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_46(11),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1915);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_8_CA_106_8x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1978,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_49(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1918);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_45_CA_69_45x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1941,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_12(45),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1881);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_17_CA_97_17x: LUT4 
  generic map(
    INIT => X"2BAF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1969,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_40(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_TEMP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1909);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_16_CA_98_16x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1970,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_41(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1910);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_13_CA_101_13x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1973,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_44(13),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1913);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_14_CA_100_14x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1972,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_43(14),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1912);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_15_CA_99_15x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1971,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_42(15),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1911);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_1_CA_113_1x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1985,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SBLSBS_1_0(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1926);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_CA_104_10x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1976,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_47(10),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1916);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_19_CA_95_19x: LUT4 
  generic map(
    INIT => X"4DDD"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_100_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1967,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_19_TRFWWBASICCELL_TEMP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1907);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_18_CA_96_18x: LUT4 
  generic map(
    INIT => X"2BAF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1968,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN31_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_39(18),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_18_TRFWWBASICCELL_TEMP2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1908);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_26_CA_88_26x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1960,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_31(26),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1900);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_32_CA_82_32x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1954,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_25(32),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1894);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_37_CA_77_37x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1949,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_20(37),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1889);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_39_CA_75_39x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1947,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_18(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1887);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_49_CA_65_49x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1937,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_8(49),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1877);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_15_0_0: MUXF6 port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_353,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_360,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(50),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_361);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_feedback_0_4x: LUT4 
  generic map(
    INIT => X"8F80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CHECKOVANDDENORM_UN20_NOTPOSSIBLEOV_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_CHECKOVANDDENORM_UN20_NOTPOSSIBLEOV_5,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN18_FEEDBACK,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_stkgen_1: LUT4_L 
  generic map(
    INIT => X"8100"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SALSBS(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN22_NOTPROP,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_1(0),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_STKGEN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un38_gen: LUT4_L 
  generic map(
    INIT => X"C080"
  )
  port map (
    I0 => N_8929,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SBLSBS(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_2(0),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SBLSBS_1(1),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN38_GEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notstickyinforsr_2: LUT4_L 
  generic map(
    INIT => X"0222"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_2_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_375x: LUT4 
  generic map(
    INIT => X"0002"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(3),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_TZ(375),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_I(375));
  x_grlfpc2_0_I_237_2: LUT4 
  generic map(
    INIT => X"0060"
  )
  port map (
    I0 => cpi_d_inst(23),
    I1 => cpi_d_inst(30),
    I2 => GRLFPC2_0_I_237_0,
    I3 => GRLFPC2_0_N_670,
    O => GRLFPC2_0_I_237_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xzCregLoadEn: LUT3 
  generic map(
    INIT => X"AB"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW86);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un1_xzybus24_s0_0_0_a2_0_0_a2: LUT3 
  generic map(
    INIT => X"10"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2354);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlbregexp_expbregloaden: LUT3 
  generic map(
    INIT => X"04"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(26),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_1(68),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_EXPBREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ctrlaregexp_exparegloaden: LUT3 
  generic map(
    INIT => X"04"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(28),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_1(68),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLOADEN);
  x_grlfpc2_0_comb_un1_rs2v: LUT4 
  generic map(
    INIT => X"4500"
  )
  port map (
    I0 => GRLFPC2_0_N_653,
    I1 => GRLFPC2_0_N_757,
    I2 => GRLFPC2_0_COMB_FPDECODE_AFQ12,
    I3 => GRLFPC2_0_COMB_RS2_1(0),
    O => GRLFPC2_0_N_750);
  x_grlfpc2_0_comb_ccwr4: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_COMB_CCWR4_1,
    I1 => GRLFPC2_0_COMB_ISFPOP2_1,
    O => GRLFPC2_0_COMB_CCWR4);
  x_grlfpc2_0_comb_lockgen_lockis2: LUT4 
  generic map(
    INIT => X"A0B0"
  )
  port map (
    I0 => GRLFPC2_0_N_776,
    I1 => GRLFPC2_0_COMB_FPDECODE_ST,
    I2 => GRLFPC2_0_COMB_LOCKGEN_LOCKI_SN_N_10,
    I3 => GRLFPC2_0_RS2_0_SQMUXA,
    O => GRLFPC2_0_N_737);
  x_grlfpc2_0_comb_un6_rs2v: LUT4 
  generic map(
    INIT => X"0045"
  )
  port map (
    I0 => GRLFPC2_0_N_653,
    I1 => GRLFPC2_0_N_757,
    I2 => GRLFPC2_0_COMB_FPDECODE_AFQ12,
    I3 => GRLFPC2_0_COMB_RS2_1(0),
    O => GRLFPC2_0_N_749);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_14_m_142x: LUT4 
  generic map(
    INIT => X"88C8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_UN17_INFORCREGSN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(144),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14_M(142));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_c_pxs_multiplexormulxff_result_0_0_2x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => N_2458,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT0(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_mixoin_1_0_0x: LUT4 
  generic map(
    INIT => X"AB01"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1869,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN22_GEN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN30_GEN,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_1(0));
  x_grlfpc2_0_comb_wrres4: LUT3 
  generic map(
    INIT => X"02"
  )
  port map (
    I0 => GRLFPC2_0_COMB_CCWR4_1,
    I1 => GRLFPC2_0_COMB_ISFPOP2_1,
    I2 => GRLFPC2_0_R_X_LD,
    O => GRLFPC2_0_COMB_WRRES4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_45: LUT4 
  generic map(
    INIT => X"8000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_39_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_43_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_41,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_45);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_46: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_39,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_40,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_46);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_47: LUT4 
  generic map(
    INIT => X"8000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_13,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_14,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_15,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_16,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_47);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_49: LUT4 
  generic map(
    INIT => X"8000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_21,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_22,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_23,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_24,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_49);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0x: LUT4 
  generic map(
    INIT => X"10D0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_853,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_854,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(57),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_4(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_2x: LUT4 
  generic map(
    INIT => X"10D0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_853,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_854,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_4(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_3x: LUT4 
  generic map(
    INIT => X"10D0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_853,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_854,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(54),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_4(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_notprop_2: LUT4 
  generic map(
    INIT => X"6006"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SBLSBS(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_2(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_2_I(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SBLSBS_1(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1809);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_gen_2: LUT3_L 
  generic map(
    INIT => X"45"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN38_GEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_2_I(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SBLSBS_1(1),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1808);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_58: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1871,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_60);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_0: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_2: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_1x: LUT4 
  generic map(
    INIT => X"10D0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_853,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_854,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(56),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_4(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_pxs_multiplexormulxff_result_0_0_am_5x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => N_2461,
    I1 => cpi_d_inst(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_71,
    O => N_12332);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_pxs_multiplexormulxff_result_0_0_bm_5x: LUT2 
  generic map(
    INIT => X"E"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTRESETORUNIMP,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(79),
    O => N_12333);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_pxs_multiplexormulxff_result_0_0_5x: MUXF5 port map (
      I0 => N_12332,
      I1 => N_12333,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1646,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_pxs_multiplexormulxff_result_0_0_am_6x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => N_2462,
    I1 => cpi_d_inst(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_71,
    O => N_12334);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_pxs_multiplexormulxff_result_0_0_bm_6x: LUT3 
  generic map(
    INIT => X"FB"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTRESETORUNIMP,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(79),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(83),
    O => N_12335);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_pxs_multiplexormulxff_result_0_0_6x: MUXF5 port map (
      I0 => N_12334,
      I1 => N_12335,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1646,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_pxs_multiplexormulxff_result_0_0_am_7x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => N_2463,
    I1 => cpi_d_inst(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_71,
    O => N_12336);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_pxs_multiplexormulxff_result_0_0_bm_7x: LUT2 
  generic map(
    INIT => X"E"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTRESETORUNIMP,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(84),
    O => N_12337);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_pxs_multiplexormulxff_result_0_0_7x: MUXF5 port map (
      I0 => N_12336,
      I1 => N_12337,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1646,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_pxs_multiplexormulxff_result_0_2_am_4x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => N_2460,
    I1 => cpi_d_inst(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_71,
    O => N_12338);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_pxs_multiplexormulxff_result_0_2_bm_4x: LUT3 
  generic map(
    INIT => X"FE"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTRESETORUNIMP,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(79),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(84),
    O => N_12339);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_pxs_multiplexormulxff_result_0_2_4x: MUXF5 port map (
      I0 => N_12338,
      I1 => N_12339,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1646,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_pxs_multiplexormulxff_result_0_2_am_2x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => N_2458,
    I1 => cpi_d_inst(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_71,
    O => N_12340);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_pxs_multiplexormulxff_result_0_2_bm_2x: LUT3 
  generic map(
    INIT => X"CD"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_OPREXCSHFT_UN3_OPREXC,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTRESETORUNIMP,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN42_CONDITIONAL,
    O => N_12341);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_pxs_multiplexormulxff_result_0_2_2x: MUXF5 port map (
      I0 => N_12340,
      I1 => N_12341,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1646,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_pxs_multiplexormulxff_result_0_2_am_1x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => N_2457,
    I1 => cpi_d_inst(9),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_71,
    O => N_12342);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_pxs_multiplexormulxff_result_0_2_bm_1x: LUT3 
  generic map(
    INIT => X"EF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTRESETORUNIMP,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN42_CONDITIONAL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1(4),
    O => N_12343);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_pxs_multiplexormulxff_result_0_2_1x: MUXF5 port map (
      I0 => N_12342,
      I1 => N_12343,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1646,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_pxs_multiplexormulxff_result_0_2_am_0x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => N_2456,
    I1 => cpi_d_inst(10),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_71,
    O => N_12344);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_pxs_multiplexormulxff_result_0_2_bm_0x: LUT4 
  generic map(
    INIT => X"CFDF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2002,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTRESETORUNIMP,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1(3),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1(4),
    O => N_12345);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_pxs_multiplexormulxff_result_0_2_0x: MUXF5 port map (
      I0 => N_12344,
      I1 => N_12345,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1646,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_89: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1901,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_89(24),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_147(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_94: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1883,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_129_1(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_129(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_96: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1884,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_130_1(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_130(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_98: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1903,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_149_1(20),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_149(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_61: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1889,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_135_1(34),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_135(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_62: LUT4 
  generic map(
    INIT => X"65A6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_62_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_66_1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1964,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_150(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_66: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1905,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_151_1(18),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_151(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_67: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1886,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_74(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_132(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_71: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1918,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_106(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_164(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_72: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1882,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_70(43),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_128(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_74: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1894,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_140_1(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_140(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_78: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1891,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_137_1(32),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_137(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_80: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1890,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_78(35),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_136(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_101: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1899,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_87(26),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_145(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_81: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1913,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_101(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_159(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_87: LUT4 
  generic map(
    INIT => X"69A5"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1907,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_95(18),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_18_TRFWWBASICCELL_TEMP2_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_153(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_68: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1923,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_111(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_83: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1921,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_109(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_167(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_105: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1920,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_108(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_166(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_73: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1919,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_107(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_165(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_93: LUT4 
  generic map(
    INIT => X"69A5"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1906,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_94(19),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_19_TRFWWBASICCELL_TEMP2_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_152(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_59: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1926,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_113(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SCLSBS(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_85: LUT4 
  generic map(
    INIT => X"C396"
  )
  port map (
    I0 => N_8825,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_64(49),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_CIN,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_UN443_CA_I,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_122(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_82: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1893,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_81(32),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_139(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_84: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1892,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_80(33),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_138(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_75: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1885,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_73(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_131(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_92: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1897,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_85(28),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_143(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_99: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1898,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_86(27),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_144(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_63: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1902,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_90(23),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_148(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_95: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1910,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_98(15),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_156(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_60: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1895,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_83(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_141(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_107: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1896,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_84(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_142(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_102: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1909,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_97(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_155(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_64: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1880,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_68(45),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_126(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_76: LUT4 
  generic map(
    INIT => X"C396"
  )
  port map (
    I0 => N_8863,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_67(46),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_CIN,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_UN462_CA_I,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_125(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_90: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1881,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_69(44),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_127(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_86: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1917,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_105(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_163(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_106: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1915,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_103(10),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_161(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_104: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1922,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_168_1(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_168(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_65: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1912,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_100(13),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_158(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_77: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1911,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_99(14),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_157(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_70: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1914,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_102(11),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_160(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_103: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1916,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_104(9),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_162(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_100: LUT4 
  generic map(
    INIT => X"69A5"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1908,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_154_1(15),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_TEMP2_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_154(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_79: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1887,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_75(38),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_133(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_69: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1888,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_76(37),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_134(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_88: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1900,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_88(25),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_146(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_1_4x: LUT4 
  generic map(
    INIT => X"9669"
  )
  port map (
    I0 => N_2362,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1872,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2122_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_1_0(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_1(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_91: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1877,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_65(48),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_123(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_97: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1878,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_66(47),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_124(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_56_si_121_48x: LUT4 
  generic map(
    INIT => X"6996"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1875,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1934,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_121_0(48),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_121(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_114: LUT4 
  generic map(
    INIT => X"6996"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_114_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1873,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1932,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2119);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_SCLSBs_1_1x: LUT4 
  generic map(
    INIT => X"6996"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_15,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1924,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1983,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SCLSBS_1(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_127x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(127),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(127));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_iv_i_a2_120x: LUT4 
  generic map(
    INIT => X"A820"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2354,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(53),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(53),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2302);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_iv_i_a2_125x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(125),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2319);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un1_xzybus24_s1_0_0_a2_0_a2: LUT4 
  generic map(
    INIT => X"0200"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un1_xzybus24_s0_0_0_a2_1_a2: LUT4 
  generic map(
    INIT => X"0100"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_173x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(173),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(173));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_118x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(118),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(118));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_iv_i_a2_116x: LUT4 
  generic map(
    INIT => X"A820"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2354,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(57),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(57),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2299);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_135x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(135),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(135));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_133x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(133),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(133));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_136x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(136),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(136));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_149x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(149),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(149));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_iv_i_a2_0_148x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(148),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2207);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_158x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(158),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(158));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_156x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(156),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(156));
  x_grlfpc2_0_v_fsr_aexc_1_sqmuxa: LUT3 
  generic map(
    INIT => X"04"
  )
  port map (
    I0 => GRLFPC2_0_COMB_CCWR4,
    I1 => GRLFPC2_0_V_FSR_AEXC_1_SQMUXA_SN,
    I2 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
    O => GRLFPC2_0_V_FSR_AEXC_1_SQMUXA);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_iv_i_a2_7_141x: LUT4 
  generic map(
    INIT => X"4000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2371);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_14_m_1_0_a2_171x: LUT4 
  generic map(
    INIT => X"0040"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14_M_1(171));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_iv_i_a2_161x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(161),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2338);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_iv_i_a2_145x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(145),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2334);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_iv_i_a2_139x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(139),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2323);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_iv_i_a2_124x: LUT4 
  generic map(
    INIT => X"A820"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2354,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(49),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(49),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2316);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_iv_i_a2_123x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(123),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2312);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_iv_i_a2_122x: LUT4 
  generic map(
    INIT => X"A820"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2354,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(51),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(51),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2309);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_iv_i_a2_121x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(121),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2305);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_rndmodeselect_un20_u_rdn: LUT4 
  generic map(
    INIT => X"000B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(21),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(1),
    I3 => GRLFPC2_0_R_FSR_RD(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN20_U_RDN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_rndmodeselect_u_rdn_1_1x: LUT4_L 
  generic map(
    INIT => X"1011"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN1_TEMP,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(2),
    I3 => GRLFPC2_0_R_FSR_RD(1),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1748);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_117x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(117),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(117));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_119x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(119),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(119));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_126x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(126),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(126));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_128x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(128),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(128));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_129x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(129),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(129));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_130x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(130),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(130));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_131x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(131),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(131));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_132x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(132),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(132));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_134x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(134),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(134));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_137x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(137),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(137));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_138x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(138),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(138));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_140x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(140),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(140));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_143x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(143),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(143));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_144x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(144),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(144));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_146x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(146),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(146));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_147x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(147),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(147));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_150x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(150),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(150));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_151x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(151),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(151));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_152x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(152),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(152));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_153x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(153),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(153));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_154x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(154),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(154));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_155x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(155),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(155));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_157x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(157),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(157));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_159x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(159),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(159));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_160x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(160),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(160));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_162x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(162),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(162));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_163x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(163),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(163));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_164x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(164),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(164));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_165x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(165),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(165));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_166x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(166),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(166));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_167x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(167),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(167));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_168x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(168),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(168));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_169x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(169),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(169));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_0_170x: LUT4 
  generic map(
    INIT => X"888C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(170),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M_0(170));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_ExpAregLoadEn: LUT4 
  generic map(
    INIT => X"FFAB"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(27),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(28),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL_1(68),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1746);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_9x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(48),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_12x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(45),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_13x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(44),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(52),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_14x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(43),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_15x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(50),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_17x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(48),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_18x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(47),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_19x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(38),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(46),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_20x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(37),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(45),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_21x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(36),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(44),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_22x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(35),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(43),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_23x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(34),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(42),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_26x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(31),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(39),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_27x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(38),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_28x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(37),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_29x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(28),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_30x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(27),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(35),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_31x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(26),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(34),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_34x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(31),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_35x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(22),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(30),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_36x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(29),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_37x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(20),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(28),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_38x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(27),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_39x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(18),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(26),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_40x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(25),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_41x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(24),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_42x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(15),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_43x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(14),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(22),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_44x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(13),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_46x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(11),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_47x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(10),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(18),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_48x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(9),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_49x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(16),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_50x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(15),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_51x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(14),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_55x: LUT3 
  generic map(
    INIT => X"8D"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_LIB(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_57x: LUT4 
  generic map(
    INIT => X"BB1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(44),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_c_pxs_multiplexormulxff_result_0_0_4x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => N_2460,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT0(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_11x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(46),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(54),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_10x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(47),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_16x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(41),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(49),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_8x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(49),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(57),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_25x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(32),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(40),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_24x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(33),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(41),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_33x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(24),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(32),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_32x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(25),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(33),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_45x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(20),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_53x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(12),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_8_0_52x: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(13),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_rndmodeselect_N_1749_i: LUT2 
  generic map(
    INIT => X"D"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN1_TEMP,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1749_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_51: LUT4_L 
  generic map(
    INIT => X"4000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_57_I_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_29,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_31,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_32,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_51);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_54: LUT4 
  generic map(
    INIT => X"4000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_56_I_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_43,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_45,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_54);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_busymulxff_un2_temp_3: LUT4 
  generic map(
    INIT => X"00A2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_BUSYMULXFF_UN2_TEMP_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN1_MIFROMINST_0,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_BUSYMULXFF_UN2_TEMP_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un53_gen: LUT4 
  generic map(
    INIT => X"00A8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SCLSBS(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(5),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN53_GEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un42_notprop: LUT4 
  generic map(
    INIT => X"AA56"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SCLSBS(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(5),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_sxdive(6),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN42_NOTPROP);
  x_grlfpc2_0_comb_v_fsr_fcc_1_m1_0_1x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_CCWR4,
    I1 => GRLFPC2_0_COMB_V_FSR_FCC_1_M0(1),
    I2 => GRLFPC2_0_R_I_CC(1),
    LO => GRLFPC2_0_COMB_V_FSR_FCC_1_M1(1));
  x_grlfpc2_0_comb_v_fsr_fcc_1_m1_0_0x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_CCWR4,
    I1 => GRLFPC2_0_COMB_V_FSR_FCC_1_M0(0),
    I2 => GRLFPC2_0_R_I_CC(0),
    LO => GRLFPC2_0_COMB_V_FSR_FCC_1_M1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_2_0_245x: LUT4 
  generic map(
    INIT => X"D8F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLOADEN_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(232),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(245),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(26),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_415);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_si_114_1_56x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1871,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_58_1(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_114_1(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_1_3x: LUT4 
  generic map(
    INIT => X"6996"
  )
  port map (
    I0 => N_2362,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_60,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2122_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_117(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_3_57x: LUT4 
  generic map(
    INIT => X"40C8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1869,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_1(57),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_STKGEN_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_3(57));
  x_grlfpc2_0_N_748_i: LUT4 
  generic map(
    INIT => X"FFBA"
  )
  port map (
    I0 => cpi_dbg_enable,
    I1 => GRLFPC2_0_N_752,
    I2 => GRLFPC2_0_COMB_RS1V_1,
    I3 => GRLFPC2_0_R_A_RF2REN(1),
    O => rfi2_ren1);
  x_grlfpc2_0_N_747_i: LUT4 
  generic map(
    INIT => X"FFBA"
  )
  port map (
    I0 => cpi_dbg_enable,
    I1 => GRLFPC2_0_N_751,
    I2 => GRLFPC2_0_COMB_RS1V_1,
    I3 => GRLFPC2_0_R_A_RF1REN(1),
    O => rfi1_ren1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_rightshifterbl_notstickyinforsr_u: LUT4 
  generic map(
    INIT => X"2023"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(42),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR);
  x_grlfpc2_0_v_fsr_aexc_2_sqmuxa: LUT4 
  generic map(
    INIT => X"0001"
  )
  port map (
    I0 => GRLFPC2_0_COMB_CCWR4,
    I1 => GRLFPC2_0_COMB_WRRES4,
    I2 => GRLFPC2_0_V_FSR_AEXC_1_SQMUXA_SN,
    I3 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
    O => GRLFPC2_0_V_FSR_AEXC_2_SQMUXA);
  x_grlfpc2_0_v_fsr_cexc_2_sqmuxa: LUT4 
  generic map(
    INIT => X"0010"
  )
  port map (
    I0 => GRLFPC2_0_COMB_CCWR4,
    I1 => GRLFPC2_0_COMB_V_I_V6,
    I2 => GRLFPC2_0_V_FSR_AEXC_1_SQMUXA_SN,
    I3 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
    O => GRLFPC2_0_V_FSR_CEXC_2_SQMUXA);
  x_grlfpc2_0_v_i_v_3_sqmuxa_272: LUT3 
  generic map(
    INIT => X"01"
  )
  port map (
    I0 => GRLFPC2_0_COMB_CCWR4,
    I1 => GRLFPC2_0_COMB_V_I_V6,
    I2 => GRLFPC2_0_COMB_WRRES4,
    O => GRLFPC2_0_N_797);
  x_grlfpc2_0_v_fsr_cexc_0_sqmuxa: LUT3 
  generic map(
    INIT => X"0E"
  )
  port map (
    I0 => GRLFPC2_0_COMB_CCWR4,
    I1 => GRLFPC2_0_COMB_WRRES4,
    I2 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
    O => GRLFPC2_0_V_FSR_CEXC_0_SQMUXA);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_iv_i_a2_172x: LUT3 
  generic map(
    INIT => X"90"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2276,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2281_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14_M_1(171),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2342);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_5x: LUT4 
  generic map(
    INIT => X"3210"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(52),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_mixoin_2_0_0x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1808,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1809,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_1(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_2(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_4x: LUT4 
  generic map(
    INIT => X"3210"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(57),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_6x: LUT4 
  generic map(
    INIT => X"3210"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_sctrl_new_10_10x: LUT4 
  generic map(
    INIT => X"4515"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN1_U_SNNOTDB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN4_TOGGLESIG,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN12_U_SNNOTDB_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1741);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_stkgen_2: LUT4_L 
  generic map(
    INIT => X"8100"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SBLSBS(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN35_NOTPROP,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_2(0),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_1(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_STKGEN_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_56: LUT4_L 
  generic map(
    INIT => X"8000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_35,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_36,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_49,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_51,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_56);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0x: LUT4 
  generic map(
    INIT => X"0100"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(57),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_1x: LUT4 
  generic map(
    INIT => X"0100"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_54_CA_117_54x: LUT4 
  generic map(
    INIT => X"B22B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1871,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_CIN_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_CIN,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_58_1(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1811);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_55_CA_116_55x: LUT4 
  generic map(
    INIT => X"B22B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1871,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_CIN,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_58_1(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1810);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_41_CA_130_41x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1884,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_130_1(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1824);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_42_CA_129_42x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1883,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_129_1(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1823);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_45_CA_126_45x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1880,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_68(45),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1820);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_51_CA_120_51x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1874,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_62(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1814);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_23_CA_148_23x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1902,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_90(23),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1842);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_25_CA_146_25x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1900,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_88(25),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1840);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_31_CA_140_31x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1894,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_140_1(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1834);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_32_CA_139_32x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1893,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_81(32),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1833);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_34_CA_137_34x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1891,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_137_1(32),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1831);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_35_CA_136_35x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1890,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_78(35),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1830);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_19_CA_152_19x: LUT4 
  generic map(
    INIT => X"2BAF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1906,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_94(19),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_19_TRFWWBASICCELL_TEMP2_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1846);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_20_CA_151_20x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1905,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_151_1(18),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1845);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_21_CA_150_21x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1904,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_150_1(19),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1844);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_temp_1x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1926,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_113(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_I(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_3_CA_168_3x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1922,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_168_1(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1862);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_49_CA_122_49x: LUT4 
  generic map(
    INIT => X"0317"
  )
  port map (
    I0 => N_8825,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_64(49),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_CIN,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_UN443_CA_I,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1816);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_50_CA_121_50x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1875,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_63(50),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1815);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_12_CA_159_12x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1913,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_101(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1853);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_26_CA_145_26x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1899,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_87(26),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1839);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_6_CA_165_6x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1919,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_107(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1859);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_5_CA_166_5x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1920,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_108(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1860);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_4_CA_167_4x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1921,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_109(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1861);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_18_CA_153_18x: LUT4 
  generic map(
    INIT => X"2BAF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1907,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_95(18),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_18_TRFWWBASICCELL_TEMP2_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1847);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_40_CA_131_40x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1885,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_73(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1825);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_39_CA_132_39x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1886,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_74(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1826);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_33_CA_138_33x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1892,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_80(33),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1832);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_30_CA_141_30x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1895,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_83(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1835);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_1_CA_170_1x: LUT4 
  generic map(
    INIT => X"48DE"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_15,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1924,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1983,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1865);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_22_CA_149_22x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1903,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_149_1(20),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1843);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_27_CA_144_27x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1898,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_86(27),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1838);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_28_CA_143_28x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1897,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_85(28),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1837);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_43_CA_128_43x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1882,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_70(43),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1822);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_29_CA_142_29x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1896,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_84(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1836);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_53_CA_118_53x: LUT4 
  generic map(
    INIT => X"B22B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1872,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_CIN_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_58_1(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1812);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_8_CA_163_8x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1917,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_105(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1857);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_10_CA_161_10x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1915,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_103(10),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1855);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_7_CA_164_7x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1918,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_106(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1858);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_46_CA_125_46x: LUT4 
  generic map(
    INIT => X"0317"
  )
  port map (
    I0 => N_8863,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_67(46),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_CIN,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_UN462_CA_I,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1819);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_44_CA_127_44x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1881,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_69(44),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1821);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_15_CA_156_15x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1910,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_98(15),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1850);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_13_CA_158_13x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1912,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_100(13),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1852);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_16_CA_155_16x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1909,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_97(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1849);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_14_CA_157_14x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1911,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_99(14),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1851);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_2_CA_169_2x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1923,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_111(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1863);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_11_CA_160_11x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1914,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_102(11),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1854);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_9_CA_162_9x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1916,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_104(9),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1856);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_17_CA_154_17x: LUT4 
  generic map(
    INIT => X"2BAF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1908,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN55_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_154_1(15),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_TEMP2_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1848);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_24_CA_147_24x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1901,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_89(24),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1841);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_36_CA_135_36x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1889,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_135_1(34),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1829);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_37_CA_134_37x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1888,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_76(37),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1828);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_38_CA_133_38x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1887,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_75(38),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1827);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_47_CA_124_47x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1878,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_66(47),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1818);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_48_CA_123_48x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1877,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_65(48),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1817);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_trfwwrray_remwtage57_52_CA_119_52x: LUT4 
  generic map(
    INIT => X"B22B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1873,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_CIN,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_58_1(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1813);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_sctrl_new_8_0_9x: LUT4 
  generic map(
    INIT => X"2F0D"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN1_TEMP,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN20_U_RDN,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(9),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_sctrl_new_8_0_8x: LUT4 
  generic map(
    INIT => X"3B31"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1748,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN1_TEMP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(8),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_42x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(38),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_48x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(44),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(48),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_am_54x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(11),
    O => N_12346);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_bm_54x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(15),
    O => N_12347);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_54x: MUXF5 port map (
      I0 => N_12346,
      I1 => N_12347,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_55x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(51),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_am_56x: LUT4 
  generic map(
    INIT => X"44E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(9),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(44),
    O => N_12348);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_bm_56x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(13),
    O => N_12349);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_56x: MUXF5 port map (
      I0 => N_12348,
      I1 => N_12349,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_57x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(53),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(57),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_8x: LUT4 
  generic map(
    INIT => X"1D11"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_44x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(40),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(44),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_52x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(48),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(52),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_50x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(46),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(50),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_46x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(42),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(46),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_40x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(36),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_20x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(16),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(20),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_18x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(14),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(18),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_17x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(13),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_15x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(11),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(15),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_14x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(10),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(14),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_13x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(9),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(13),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_12x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_11x: LUT4 
  generic map(
    INIT => X"1D11"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(11),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(50),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_4_0_10x: LUT4 
  generic map(
    INIT => X"1D11"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(10),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_NE_10: LUT4 
  generic map(
    INIT => X"0906"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_3,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_NE_10);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_2_sqmuxa: LUT4 
  generic map(
    INIT => X"5D55"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLOADEN_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(25),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(26),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA);
  x_grlfpc2_0_v_fsr_cexc_3_sqmuxa: LUT3 
  generic map(
    INIT => X"02"
  )
  port map (
    I0 => GRLFPC2_0_N_797,
    I1 => GRLFPC2_0_V_FSR_AEXC_1_SQMUXA_SN,
    I2 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
    O => GRLFPC2_0_V_FSR_CEXC_3_SQMUXA);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m3_1: LUT4 
  generic map(
    INIT => X"3313"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLOADEN_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(27),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(28),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_800);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_2x: LUT4 
  generic map(
    INIT => X"CEDF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_4(0),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_4(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_3x: LUT4 
  generic map(
    INIT => X"CEDF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_4(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_4(3),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1: LUT4 
  generic map(
    INIT => X"8000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_46,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_47,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_54,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_56,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_14_m_171x: LUT4 
  generic map(
    INIT => X"40C0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2276,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14_M_0(171),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14_M_1(171),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_T_3_I_A2_0_0(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_14_M(171));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_iv_i_a2_0_141x: LUT3 
  generic map(
    INIT => X"40"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2276,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2371,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_T_3_I_A2_0_0(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2328);
  x_grlfpc2_0_comb_wren2_9_iv: LUT4 
  generic map(
    INIT => X"10F0"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_COMB_WRADDR_5(0),
    I2 => GRLFPC2_0_COMB_WREN2_9_IV_0,
    I3 => GRLFPC2_0_COMB_WRRES4,
    O => GRLFPC2_0_N_708);
  x_grlfpc2_0_comb_wren1_9_iv_0: LUT3 
  generic map(
    INIT => X"4F"
  )
  port map (
    I0 => GRLFPC2_0_COMB_RDD_3,
    I1 => GRLFPC2_0_COMB_WRADDR_5(0),
    I2 => GRLFPC2_0_COMB_WRRES4,
    O => GRLFPC2_0_COMB_WREN1_9_IV_0);
  x_grlfpc2_0_comb_v_fsr_aexc_1_iv_0_3x: LUT4_L 
  generic map(
    INIT => X"153F"
  )
  port map (
    I0 => cpi_dbg_data(8),
    I1 => cpi_lddata(8),
    I2 => GRLFPC2_0_V_FSR_AEXC_1_SQMUXA,
    I3 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
    LO => GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_0(3));
  x_grlfpc2_0_comb_v_fsr_aexc_1_iv_0_0x: LUT4_L 
  generic map(
    INIT => X"153F"
  )
  port map (
    I0 => cpi_dbg_data(5),
    I1 => cpi_lddata(5),
    I2 => GRLFPC2_0_V_FSR_AEXC_1_SQMUXA,
    I3 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
    LO => GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_0(0));
  x_grlfpc2_0_comb_v_fsr_aexc_1_iv_0_2x: LUT4_L 
  generic map(
    INIT => X"153F"
  )
  port map (
    I0 => cpi_dbg_data(7),
    I1 => cpi_lddata(7),
    I2 => GRLFPC2_0_V_FSR_AEXC_1_SQMUXA,
    I3 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
    LO => GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_0(2));
  x_grlfpc2_0_comb_v_fsr_aexc_1_iv_0_4x: LUT4_L 
  generic map(
    INIT => X"153F"
  )
  port map (
    I0 => cpi_dbg_data(9),
    I1 => cpi_lddata(9),
    I2 => GRLFPC2_0_V_FSR_AEXC_1_SQMUXA,
    I3 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
    LO => GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_0(4));
  x_grlfpc2_0_comb_v_fsr_aexc_1_iv_0_1x: LUT4_L 
  generic map(
    INIT => X"153F"
  )
  port map (
    I0 => cpi_dbg_data(6),
    I1 => cpi_lddata(6),
    I2 => GRLFPC2_0_V_FSR_AEXC_1_SQMUXA,
    I3 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
    LO => GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_0(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_83_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(137),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(38),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_83_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_60_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(130),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(45),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_60_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_95_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(155),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(20),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_95_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_61_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(129),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(46),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_61_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_74_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(146),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(29),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_74_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_59_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(131),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(44),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_59_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_94_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(156),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(19),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_94_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_58_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(132),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(43),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_58_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_109_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(168),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(7),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_109_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_82_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(138),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(37),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_82_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_71_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(119),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(56),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_71_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_87_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(163),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(12),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_87_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_97_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(153),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(22),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_97_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_96_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(154),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(21),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_96_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_84_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(136),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(39),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_84_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_73_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(147),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(28),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_73_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_72_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(148),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(27),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_72_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_81_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(139),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(36),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_81_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_112_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(165),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(10),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_112_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_113_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(164),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(11),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_113_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_110_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(167),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(8),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_110_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_106_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(171),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(4),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_106_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_105_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(172),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(3),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_105_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_101_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(149),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(26),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_101_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_99_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(151),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(24),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_99_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_86_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(134),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(41),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_86_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_85_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(135),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(40),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_85_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_88_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(162),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(13),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_88_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_79_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(141),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(34),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_79_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_108_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(169),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(6),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_108_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_62_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(128),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(47),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_62_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_80_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(140),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(35),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_80_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_65_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(125),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(50),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_65_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_93_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(157),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(18),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_93_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_111_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(166),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(9),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_111_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_67_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(123),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(52),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_67_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_78_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(142),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(33),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_78_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_69_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(121),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(54),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_69_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_98_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(152),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(23),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_98_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_75_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(145),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(30),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_75_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_70_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(120),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(55),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_70_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_90_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(160),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(15),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_90_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_57_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(133),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(42),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_57_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_63_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(127),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(48),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_63_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_89_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(161),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(14),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_89_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_91_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(159),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(16),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_91_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_107_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(170),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(5),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_107_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_92_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(158),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(17),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_92_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_103_0: LUT4_L 
  generic map(
    INIT => X"57DF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2354,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(1),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_103_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_76_0: LUT4_L 
  generic map(
    INIT => X"57DF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2354,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(31),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(31),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_76_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_104_0: LUT4_L 
  generic map(
    INIT => X"57DF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2354,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(2),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(2),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_104_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_77_0: LUT4_L 
  generic map(
    INIT => X"5515"
  )
  port map (
    I0 => N_2376,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(143),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_77_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_77_1: LUT4 
  generic map(
    INIT => X"57DF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2354,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(32),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(32),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_77_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_4x: LUT4 
  generic map(
    INIT => X"D1DD"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(4),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_4(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_5x: LUT4 
  generic map(
    INIT => X"D1DD"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(5),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_4(3),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_6x: LUT4 
  generic map(
    INIT => X"CDEF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    O => N_12350);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_6x: LUT4 
  generic map(
    INIT => X"CDEF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(57),
    O => N_12351);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_6x: MUXF5 port map (
      I0 => N_12350,
      I1 => N_12351,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_7x: LUT4 
  generic map(
    INIT => X"CDEF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(50),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(54),
    O => N_12352);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_7x: LUT4 
  generic map(
    INIT => X"CDEF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(52),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(56),
    O => N_12353);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_7x: MUXF5 port map (
      I0 => N_12352,
      I1 => N_12353,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un49_notprop: LUT4 
  generic map(
    INIT => X"399C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1926,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SCLSBS_1(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_CIN_3,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_113(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN49_NOTPROP);
  x_grlfpc2_0_r_mk_ldopc_1: LUT4 
  generic map(
    INIT => X"4051"
  )
  port map (
    I0 => CPO_EXC_INT_2,
    I1 => GRLFPC2_0_N_737,
    I2 => GRLFPC2_0_N_777,
    I3 => GRLFPC2_0_COMB_LOCKGEN_LOCKI_SN_N_10,
    O => GRLFPC2_0_R_MK_LDOPC_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_49_1_258x: LUT4 
  generic map(
    INIT => X"9669"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1810,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1871,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1932,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_49_1_2(258),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_49_1(258));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_31x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1840,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_145(24),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_26x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1835,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_140(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_55x: LUT4 
  generic map(
    INIT => X"6A95"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1865,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_TEMP2_3,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_52x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1861,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_166(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_51x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1860,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_165(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_50x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1859,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_164(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_47x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1856,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_161(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_46x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1855,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_160(9),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_44x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1853,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_158(11),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_41x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1850,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_155(14),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_25x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1834,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_139(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_23x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1832,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_137(32),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_22x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1831,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_136(33),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_21x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1830,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_135(34),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_19x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1828,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_133(36),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_18x: LUT4 
  generic map(
    INIT => X"69A5"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1827,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_132(37),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_TEMP2_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_16x: LUT4 
  generic map(
    INIT => X"69A5"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1825,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_130(39),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_TEMP2_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_15x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1824,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_129(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_14x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1823,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_128(41),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_11x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1820,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_125(44),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_37x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1846,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_151(18),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_18_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_36x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1845,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_150(19),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_19_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_35x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1844,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_149(20),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_33x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1842,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_147(22),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_7x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1816,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_121(48),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_NE: LUT4 
  generic map(
    INIT => X"1000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_NE_7,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_NE_10,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_8x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1817,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_122(47),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(8));
  x_grlfpc2_0_comb_lock_1: LUT4 
  generic map(
    INIT => X"7020"
  )
  port map (
    I0 => GRLFPC2_0_N_737,
    I1 => GRLFPC2_0_N_777,
    I2 => GRLFPC2_0_COMB_LOCK_1_1_0,
    I3 => GRLFPC2_0_COMB_LOCKGEN_LOCKI_SN_N_10,
    O => cpo_ldlock);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_45x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1854,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_159(10),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_29x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1838,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_143(26),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_17x: LUT4 
  generic map(
    INIT => X"69A5"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1826,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_131(38),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_TEMP2_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_38x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1847,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_152(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_10x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1819,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_124(45),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_24x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1833,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_138(31),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_30x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1839,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_144(25),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_34x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1843,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_148(21),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_42x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1851,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_156(13),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_49x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1858,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_163(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_27x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1836,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_141(28),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_28x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1837,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_142(27),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_13x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1822,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_127(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_43x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1852,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_157(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_12x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1821,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_126(43),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_53x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1862,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_167(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_54x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1863,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_168(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_48x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1857,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_162(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_40x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1849,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_154(15),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_39x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1848,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_153(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_20x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1829,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_134(35),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_32x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1841,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_146(23),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_3x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1812,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_117(52),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_4x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1813,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_1(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_6x: LUT4 
  generic map(
    INIT => X"6996"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1815,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1874,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_120_1(49),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_9x: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1818,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_123(46),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_2x: LUT4 
  generic map(
    INIT => X"9669"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1811,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_CIN,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_114_1(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_5x: LUT4 
  generic map(
    INIT => X"9669"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1814,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2119,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_CIN_2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_114_1_1_0(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(5));
  x_grlfpc2_0_v_i_v_3_sqmuxa_i: LUT3 
  generic map(
    INIT => X"7F"
  )
  port map (
    I0 => GRLFPC2_0_N_762,
    I1 => GRLFPC2_0_N_797,
    I2 => GRLFPC2_0_V_I_EXEC26,
    O => GRLFPC2_0_V_I_V_3_SQMUXA_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m3: LUT4 
  generic map(
    INIT => X"A22A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLOADEN_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(25),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(26),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m5: LUT4 
  generic map(
    INIT => X"0507"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1746,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(27),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_815);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_9x: LUT4 
  generic map(
    INIT => X"E2EE"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(9),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(52),
    O => N_12354);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_9x: LUT4 
  generic map(
    INIT => X"CDEF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(50),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(54),
    O => N_12355);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_9x: MUXF5 port map (
      I0 => N_12354,
      I1 => N_12355,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_10x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(10),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_11x: LUT4 
  generic map(
    INIT => X"E2EE"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(11),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(50),
    O => N_12356);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_11x: LUT4 
  generic map(
    INIT => X"E2EE"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(9),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(52),
    O => N_12357);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_11x: MUXF5 port map (
      I0 => N_12356,
      I1 => N_12357,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_13x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(11),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(13),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_15x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(13),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(15),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_16x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(12),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12358);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_16x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(10),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(14),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12359);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_16x: MUXF5 port map (
      I0 => N_12358,
      I1 => N_12359,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_17x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(15),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_18x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(14),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(18),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12360);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_18x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(12),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12361);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_18x: MUXF5 port map (
      I0 => N_12360,
      I1 => N_12361,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_19x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(15),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(19),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12362);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_19x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(13),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12363);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_19x: MUXF5 port map (
      I0 => N_12362,
      I1 => N_12363,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_21x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(17),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(21),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12364);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_21x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(15),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(19),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12365);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_21x: MUXF5 port map (
      I0 => N_12364,
      I1 => N_12365,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_22x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(18),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(22),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12366);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_22x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(16),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(20),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12367);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_22x: MUXF5 port map (
      I0 => N_12366,
      I1 => N_12367,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_23x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(19),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(23),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12368);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_23x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(17),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(21),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12369);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_23x: MUXF5 port map (
      I0 => N_12368,
      I1 => N_12369,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_24x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(20),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(24),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12370);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_24x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(18),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(22),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12371);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_24x: MUXF5 port map (
      I0 => N_12370,
      I1 => N_12371,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_25x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(25),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12372);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_25x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(19),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(23),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12373);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_25x: MUXF5 port map (
      I0 => N_12372,
      I1 => N_12373,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_26x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(22),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(26),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12374);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_26x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(20),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(24),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12375);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_26x: MUXF5 port map (
      I0 => N_12374,
      I1 => N_12375,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_27x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(27),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12376);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_27x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(25),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12377);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_27x: MUXF5 port map (
      I0 => N_12376,
      I1 => N_12377,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_28x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(24),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(28),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12378);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_28x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(22),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(26),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12379);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_28x: MUXF5 port map (
      I0 => N_12378,
      I1 => N_12379,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_29x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(25),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12380);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_29x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(27),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12381);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_29x: MUXF5 port map (
      I0 => N_12380,
      I1 => N_12381,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_30x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(26),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12382);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_30x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(24),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(28),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12383);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_30x: MUXF5 port map (
      I0 => N_12382,
      I1 => N_12383,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_31x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(27),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(31),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12384);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_31x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(25),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12385);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_31x: MUXF5 port map (
      I0 => N_12384,
      I1 => N_12385,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_32x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(28),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(32),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12386);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_32x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(26),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12387);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_32x: MUXF5 port map (
      I0 => N_12386,
      I1 => N_12387,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_33x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(29),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(33),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12388);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_33x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(27),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(31),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12389);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_33x: MUXF5 port map (
      I0 => N_12388,
      I1 => N_12389,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_34x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(34),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12390);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_34x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(28),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(32),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12391);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_34x: MUXF5 port map (
      I0 => N_12390,
      I1 => N_12391,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_35x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(31),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(35),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12392);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_35x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(29),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(33),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12393);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_35x: MUXF5 port map (
      I0 => N_12392,
      I1 => N_12393,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_36x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(32),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(36),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12394);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_36x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(34),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12395);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_36x: MUXF5 port map (
      I0 => N_12394,
      I1 => N_12395,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_37x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(33),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(37),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12396);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_37x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(31),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(35),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12397);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_37x: MUXF5 port map (
      I0 => N_12396,
      I1 => N_12397,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_38x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(34),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(38),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12398);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_38x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(32),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(36),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12399);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_38x: MUXF5 port map (
      I0 => N_12398,
      I1 => N_12399,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_39x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(35),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12400);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_39x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(33),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(37),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12401);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_39x: MUXF5 port map (
      I0 => N_12400,
      I1 => N_12401,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_40x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(36),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12402);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_40x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(34),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(38),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12403);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_40x: MUXF5 port map (
      I0 => N_12402,
      I1 => N_12403,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_41x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(37),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(41),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12404);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_41x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(35),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12405);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_41x: MUXF5 port map (
      I0 => N_12404,
      I1 => N_12405,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_43x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(39),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(43),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12406);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_43x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(37),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(41),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12407);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_43x: MUXF5 port map (
      I0 => N_12406,
      I1 => N_12407,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_45x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(41),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(45),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12408);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_45x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(39),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(43),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12409);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_45x: MUXF5 port map (
      I0 => N_12408,
      I1 => N_12409,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_46x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(44),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(46),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_47x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(43),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(47),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12410);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_47x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(41),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(45),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12411);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_47x: MUXF5 port map (
      I0 => N_12410,
      I1 => N_12411,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_49x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(45),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(49),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12412);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_49x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(43),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(47),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12413);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_49x: MUXF5 port map (
      I0 => N_12412,
      I1 => N_12413,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_51x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(47),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12414);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_51x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(45),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(49),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12415);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_51x: MUXF5 port map (
      I0 => N_12414,
      I1 => N_12415,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_53x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(49),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12416);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_53x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(47),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12417);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_53x: MUXF5 port map (
      I0 => N_12416,
      I1 => N_12417,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_54x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(52),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(54),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_am_55x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(51),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12418);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_bm_55x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(49),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_8(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    O => N_12419);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_55x: MUXF5 port map (
      I0 => N_12418,
      I1 => N_12419,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_56x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(54),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(56),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_52x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(50),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(52),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_50x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(48),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(50),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_48x: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(46),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(48),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(48));
  x_grlfpc2_0_comb_v_fsr_aexc_1_iv_1_3x: LUT3_L 
  generic map(
    INIT => X"2A"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_0(3),
    I1 => GRLFPC2_0_R_FSR_AEXC(3),
    I2 => GRLFPC2_0_V_FSR_AEXC_2_SQMUXA,
    LO => GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_1(3));
  x_grlfpc2_0_comb_v_fsr_aexc_1_iv_1_0x: LUT3_L 
  generic map(
    INIT => X"2A"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_0(0),
    I1 => GRLFPC2_0_R_FSR_AEXC(0),
    I2 => GRLFPC2_0_V_FSR_AEXC_2_SQMUXA,
    LO => GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_1(0));
  x_grlfpc2_0_comb_v_fsr_aexc_1_iv_1_2x: LUT3_L 
  generic map(
    INIT => X"2A"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_0(2),
    I1 => GRLFPC2_0_R_FSR_AEXC(2),
    I2 => GRLFPC2_0_V_FSR_AEXC_2_SQMUXA,
    LO => GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_1(2));
  x_grlfpc2_0_comb_v_fsr_aexc_1_iv_1_4x: LUT3_L 
  generic map(
    INIT => X"2A"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_0(4),
    I1 => GRLFPC2_0_R_FSR_AEXC(4),
    I2 => GRLFPC2_0_V_FSR_AEXC_2_SQMUXA,
    LO => GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_1(4));
  x_grlfpc2_0_comb_v_fsr_aexc_1_iv_1_1x: LUT3_L 
  generic map(
    INIT => X"2A"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_0(1),
    I1 => GRLFPC2_0_R_FSR_AEXC(1),
    I2 => GRLFPC2_0_V_FSR_AEXC_2_SQMUXA,
    LO => GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_1(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_5_57x: LUT4 
  generic map(
    INIT => X"40C8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1809,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_3(57),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_STKGEN_2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_1(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_5(57));
  x_grlfpc2_0_N_745_i: LUT4 
  generic map(
    INIT => X"FFBA"
  )
  port map (
    I0 => cpi_dbg_enable,
    I1 => GRLFPC2_0_N_749,
    I2 => GRLFPC2_0_COMB_FPDECODE_AFQ12,
    I3 => GRLFPC2_0_R_A_RF2REN(2),
    O => rfi2_ren2);
  x_grlfpc2_0_N_746_i: LUT4 
  generic map(
    INIT => X"FFBA"
  )
  port map (
    I0 => cpi_dbg_enable,
    I1 => GRLFPC2_0_N_750,
    I2 => GRLFPC2_0_COMB_FPDECODE_AFQ12,
    I3 => GRLFPC2_0_R_A_RF1REN(2),
    O => rfi1_ren2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_244x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_FPO_EXP(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_OP2(52),
    O => N_12420);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_244x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(244),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(257),
    O => N_12421);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_244x: MUXF5 port map (
      I0 => N_12420,
      I1 => N_12421,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_800,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_802);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_243x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_FPO_EXP(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_OP2(53),
    O => N_12422);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_243x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(243),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(256),
    O => N_12423);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_243x: MUXF5 port map (
      I0 => N_12422,
      I1 => N_12423,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_800,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_803);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_242x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_FPO_EXP(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_OP2(54),
    O => N_12424);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_242x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(242),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(255),
    O => N_12425);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_242x: MUXF5 port map (
      I0 => N_12424,
      I1 => N_12425,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_800,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_804);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_241x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_FPO_EXP(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_OP2(55),
    O => N_12426);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_241x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(241),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(254),
    O => N_12427);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_241x: MUXF5 port map (
      I0 => N_12426,
      I1 => N_12427,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_800,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_805);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_239x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_FPO_EXP(5),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_OP2(57),
    O => N_12428);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_239x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(239),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(252),
    O => N_12429);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_239x: MUXF5 port map (
      I0 => N_12428,
      I1 => N_12429,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_800,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_807);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_238x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_FPO_EXP(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_OP2(58),
    O => N_12430);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_238x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(238),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(251),
    O => N_12431);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_238x: MUXF5 port map (
      I0 => N_12430,
      I1 => N_12431,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_800,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_808);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_237x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_FPO_EXP(7),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_OP2(59),
    O => N_12432);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_237x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(237),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(250),
    O => N_12433);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_237x: MUXF5 port map (
      I0 => N_12432,
      I1 => N_12433,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_800,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_809);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_236x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_FPO_EXP(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_OP2(60),
    O => N_12434);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_236x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(236),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(249),
    O => N_12435);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_236x: MUXF5 port map (
      I0 => N_12434,
      I1 => N_12435,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_800,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_810);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_235x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_FPO_EXP(9),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_OP2(61),
    O => N_12436);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_235x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(235),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(248),
    O => N_12437);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_235x: MUXF5 port map (
      I0 => N_12436,
      I1 => N_12437,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_800,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_811);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_234x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_FPO_EXP(10),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_OP2(62),
    O => N_12438);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_234x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(234),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(247),
    O => N_12439);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_234x: MUXF5 port map (
      I0 => N_12438,
      I1 => N_12439,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_800,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_812);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_233x: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => N_2476,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    O => N_12440);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_233x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(233),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(246),
    O => N_12441);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_233x: MUXF5 port map (
      I0 => N_12440,
      I1 => N_12441,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_800,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_813);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_232x: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => N_2477,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    O => N_12442);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_232x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(232),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(245),
    O => N_12443);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_232x: MUXF5 port map (
      I0 => N_12442,
      I1 => N_12443,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_800,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_814);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_feedback_0_3x: LUT3 
  generic map(
    INIT => X"B8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN18_FEEDBACK,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(57),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_240x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_FPO_EXP(4),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_OP2(56),
    O => N_12444);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_240x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLAREGEXP_EXPAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(240),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(253),
    O => N_12445);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_240x: MUXF5 port map (
      I0 => N_12444,
      I1 => N_12445,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_800,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_806);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_1x: LUT2 
  generic map(
    INIT => X"6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_49_1(258),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_0x: LUT2 
  generic map(
    INIT => X"6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_49_1(258),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(0));
  x_grlfpc2_0_comb_wren1_9_iv: LUT4 
  generic map(
    INIT => X"080C"
  )
  port map (
    I0 => cpi_x_inst(25),
    I1 => GRLFPC2_0_COMB_WREN1_9_IV_0,
    I2 => GRLFPC2_0_WREN1_1_SQMUXA_1,
    I3 => GRLFPC2_0_WREN2_2_SQMUXA,
    O => GRLFPC2_0_N_707);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_gen_3: LUT3 
  generic map(
    INIT => X"4D"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN53_GEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_I(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SCLSBS_1(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1743);
  x_grlfpc2_0_comb_fpop_1: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_R_MK_LDOPC_1,
    I1 => GRLFPC2_0_R_MK_LDOPC_2,
    I2 => GRLFPC2_0_RS2_0_SQMUXA,
    O => GRLFPC2_0_COMB_FPOP_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_101x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1853,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_158(11),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1763);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_103x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1855,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_160(9),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1761);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_104x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1856,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_161(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1760);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_107x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1859,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_164(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1757);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_108x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1860,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_165(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1756);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_109x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1861,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_166(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1755);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_112x: LUT4 
  generic map(
    INIT => X"2ABF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1865,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_TEMP2_3,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1752);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_88x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1840,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_145(24),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1776);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_90x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1842,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_147(22),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1774);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_92x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1844,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_149(20),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1772);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_93x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1845,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_150(19),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_19_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1771);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_98x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1850,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_155(14),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1766);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_71x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1823,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_128(41),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1793);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_73x: LUT4 
  generic map(
    INIT => X"2BAF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1825,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_130(39),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_TEMP2_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1791);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_75x: LUT4 
  generic map(
    INIT => X"2BAF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1827,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_132(37),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_TEMP2_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1789);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_78x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1830,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_135(34),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1786);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_79x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1831,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_136(33),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1785);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_83x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1835,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_140(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1781);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_58x: LUT4 
  generic map(
    INIT => X"B22B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1810,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_CIN_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_114_1(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1806);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_59x: LUT4 
  generic map(
    INIT => X"B22B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1811,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_CIN,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_114_1(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1805);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_62x: LUT4 
  generic map(
    INIT => X"8E2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1814,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2119,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_CIN_2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_114_1_1_0(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1802);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_63x: LUT4 
  generic map(
    INIT => X"28BE"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1815,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1874,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_120_1(49),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1801);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_65x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1817,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_122(47),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1799);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_68x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1820,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_125(44),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1796);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_86x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1838,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_143(26),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1778);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_102x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1854,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_159(10),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1762);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_95x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1847,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_152(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1769);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_74x: LUT4 
  generic map(
    INIT => X"2BAF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1826,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_131(38),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_TEMP2_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1790);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_81x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1833,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_138(31),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1783);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_82x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1834,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_139(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1782);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_91x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1843,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_148(21),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1773);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_87x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1839,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_144(25),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1777);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_85x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1837,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_142(27),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1779);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_84x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1836,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_141(28),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1780);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_106x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1858,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_163(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_CIN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1758);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_69x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1821,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_126(43),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1795);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_110x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1862,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_167(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1754);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_105x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1857,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_162(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_CIN_2,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1759);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_96x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1848,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_153(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1768);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_77x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1829,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_134(35),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_CIN_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1787);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_61x: LUT3 
  generic map(
    INIT => X"2B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1813,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_1(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_CIN_3,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1803);
  x_grlfpc2_0_comb_wren2_1_0: LUT4 
  generic map(
    INIT => X"A3A0"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => GRLFPC2_0_N_708,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    I3 => holdn,
    O => rfi2_wren);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_246x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => N_2476,
    I1 => N_2477,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_EXPBREGLC_1(1),
    O => N_12446);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_246x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_EXPBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(233),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(246),
    O => N_12447);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_246x: MUXF5 port map (
      I0 => N_12446,
      I1 => N_12447,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_428);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_247x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => N_2476,
    I1 => GRLFPC2_0_FPO_EXP(10),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_EXPBREGLC_1(1),
    O => N_12448);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_247x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_EXPBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(234),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(247),
    O => N_12449);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_247x: MUXF5 port map (
      I0 => N_12448,
      I1 => N_12449,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_427);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_248x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_EXP(9),
    I1 => GRLFPC2_0_FPO_EXP(10),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_EXPBREGLC_1(1),
    O => N_12450);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_248x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_EXPBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(235),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(248),
    O => N_12451);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_248x: MUXF5 port map (
      I0 => N_12450,
      I1 => N_12451,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_426);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_249x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_EXP(8),
    I1 => GRLFPC2_0_FPO_EXP(9),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_EXPBREGLC_1(1),
    O => N_12452);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_249x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_EXPBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(236),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(249),
    O => N_12453);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_249x: MUXF5 port map (
      I0 => N_12452,
      I1 => N_12453,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_425);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_252x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_EXP(5),
    I1 => GRLFPC2_0_FPO_EXP(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_EXPBREGLC_1(1),
    O => N_12454);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_252x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_EXPBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(239),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(252),
    O => N_12455);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_252x: MUXF5 port map (
      I0 => N_12454,
      I1 => N_12455,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_422);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_254x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_EXP(3),
    I1 => GRLFPC2_0_FPO_EXP(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_EXPBREGLC_1(1),
    O => N_12456);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_254x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_EXPBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(241),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(254),
    O => N_12457);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_254x: MUXF5 port map (
      I0 => N_12456,
      I1 => N_12457,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_420);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_255x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_EXP(2),
    I1 => GRLFPC2_0_FPO_EXP(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_EXPBREGLC_1(1),
    O => N_12458);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_255x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_EXPBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(242),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(255),
    O => N_12459);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_255x: MUXF5 port map (
      I0 => N_12458,
      I1 => N_12459,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_419);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_257x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_FPO_EXP(0),
    I1 => GRLFPC2_0_FPO_EXP(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA,
    O => N_12460);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_257x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_EXPBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(244),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(257),
    O => N_12461);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_257x: MUXF5 port map (
      I0 => N_12460,
      I1 => N_12461,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_417);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_256x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_FPO_EXP(1),
    I1 => GRLFPC2_0_FPO_EXP(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA,
    O => N_12462);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_256x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_EXPBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(243),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(256),
    O => N_12463);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_256x: MUXF5 port map (
      I0 => N_12462,
      I1 => N_12463,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_418);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_253x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_FPO_EXP(4),
    I1 => GRLFPC2_0_FPO_EXP(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA,
    O => N_12464);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_253x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_EXPBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(240),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(253),
    O => N_12465);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_253x: MUXF5 port map (
      I0 => N_12464,
      I1 => N_12465,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_421);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_251x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_FPO_EXP(6),
    I1 => GRLFPC2_0_FPO_EXP(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA,
    O => N_12466);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_251x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_EXPBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(238),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(251),
    O => N_12467);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_251x: MUXF5 port map (
      I0 => N_12466,
      I1 => N_12467,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_423);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_250x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_FPO_EXP(7),
    I1 => GRLFPC2_0_FPO_EXP(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA,
    O => N_12468);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_250x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLBREGEXP_EXPBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(237),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(250),
    O => N_12469);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_250x: MUXF5 port map (
      I0 => N_12468,
      I1 => N_12469,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_424);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_feedback_0_0_1x: LUT4_L 
  generic map(
    INIT => X"FE0E"
  )
  port map (
    I0 => N_2477,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN19_FEEDBACK_2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_AREGXORBREG,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_344);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_un28_stkout: LUT4 
  generic map(
    INIT => X"3677"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN42_NOTPROP,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN49_NOTPROP,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN53_GEN,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_2(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN28_STKOUT);
  x_grlfpc2_0_fpi_start: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_N_782,
    I1 => GRLFPC2_0_COMB_FPOP_1,
    I2 => holdn,
    O => GRLFPC2_0_FPI_START);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_am_100x: LUT2 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => rfo2_data1(12),
    O => N_12470);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_bm_100x: LUT3 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1852,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_157(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_CIN,
    O => N_12471);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_100x: MUXF5 port map (
      I0 => N_12470,
      I1 => N_12471,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_459);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_am_97x: LUT2 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => rfo2_data1(15),
    O => N_12472);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_bm_97x: LUT3 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1849,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_154(15),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_CIN_3,
    O => N_12473);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_97x: MUXF5 port map (
      I0 => N_12472,
      I1 => N_12473,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_462);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_am_94x: LUT2 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => rfo2_data1(18),
    O => N_12474);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_bm_94x: LUT3 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1846,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_151(18),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_18_TRFWWBASICCELL_CIN,
    O => N_12475);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_94x: MUXF5 port map (
      I0 => N_12474,
      I1 => N_12475,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_465);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_am_80x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP1(32),
    I2 => GRLFPC2_0_OP1(35),
    O => N_12476);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_bm_80x: LUT3 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1832,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_137(32),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_CIN_2,
    O => N_12477);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_80x: MUXF5 port map (
      I0 => N_12476,
      I1 => N_12477,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_479);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_am_76x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP1(36),
    I2 => GRLFPC2_0_OP1(39),
    O => N_12478);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_bm_76x: LUT3 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1828,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_133(36),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_CIN_2,
    O => N_12479);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_76x: MUXF5 port map (
      I0 => N_12478,
      I1 => N_12479,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_483);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_am_72x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP1(40),
    I2 => GRLFPC2_0_OP1(43),
    O => N_12480);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_bm_72x: LUT3 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1824,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_129(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_CIN,
    O => N_12481);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_72x: MUXF5 port map (
      I0 => N_12480,
      I1 => N_12481,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_487);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_am_66x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP1(46),
    I2 => GRLFPC2_0_OP1(49),
    O => N_12482);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_bm_66x: LUT3 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1818,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_123(46),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_CIN_1,
    O => N_12483);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_66x: MUXF5 port map (
      I0 => N_12482,
      I1 => N_12483,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_493);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_am_64x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP1(48),
    I2 => GRLFPC2_0_OP1(51),
    O => N_12484);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_bm_64x: LUT3 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1816,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_121(48),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_CIN_3,
    O => N_12485);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_64x: MUXF5 port map (
      I0 => N_12484,
      I1 => N_12485,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_495);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_mixoin_3_0_0x: LUT4 
  generic map(
    INIT => X"EA2A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1743,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN42_NOTPROP,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN49_NOTPROP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_2(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_3(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_am_70x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP1(42),
    I2 => GRLFPC2_0_OP1(45),
    O => N_12486);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_bm_70x: LUT3 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1822,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_127(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_CIN_2,
    O => N_12487);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_70x: MUXF5 port map (
      I0 => N_12486,
      I1 => N_12487,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_489);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_am_111x: LUT2 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => rfo2_data1(1),
    O => N_12488);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_bm_111x: LUT3 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1863,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_168(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_CIN_1,
    O => N_12489);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_111x: MUXF5 port map (
      I0 => N_12488,
      I1 => N_12489,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_448);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_am_67x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => GRLFPC2_0_OP1(45),
    I2 => GRLFPC2_0_OP1(48),
    O => N_12490);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_bm_67x: LUT3 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1819,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_124(45),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_CIN_1,
    O => N_12491);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_67x: MUXF5 port map (
      I0 => N_12490,
      I1 => N_12491,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_492);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_am_99x: LUT2 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => rfo2_data1(13),
    O => N_12492);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_bm_99x: LUT3 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1851,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_156(13),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_CIN_1,
    O => N_12493);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_99x: MUXF5 port map (
      I0 => N_12492,
      I1 => N_12493,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_460);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_am_89x: LUT2 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I1 => rfo2_data1(23),
    O => N_12494);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_bm_89x: LUT3 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1841,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_146(23),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_CIN_3,
    O => N_12495);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_89x: MUXF5 port map (
      I0 => N_12494,
      I1 => N_12495,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_470);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_r_sctrl_3_sn_m4_0: LUT3 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_I(22),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1529);
  x_grlfpc2_0_comb_wren1_1_0: LUT4 
  generic map(
    INIT => X"5350"
  )
  port map (
    I0 => cpi_dbg_addr(0),
    I1 => GRLFPC2_0_N_707,
    I2 => GRLFPC2_0_WRADDR_0_SQMUXA,
    I3 => holdn,
    O => rfi1_wren);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_feedback_u_0_1x: LUT4 
  generic map(
    INIT => X"ABA8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_344,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN18_FEEDBACK,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN19_FEEDBACK,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(59),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_57x: LUT4 
  generic map(
    INIT => X"0222"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_5(57),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN28_STKOUT,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN42_NOTPROP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_2(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1724);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_m_3x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_M(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_4x: LUT3 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2023,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_m_6x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_M(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_m_9x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(9),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_M(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_19x: LUT3 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2023,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_m_20x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(20),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_M(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_54x: LUT3 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2023,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(54),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m4_0: LUT4 
  generic map(
    INIT => X"2AAA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA_M1_E_0,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(5),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_5x: LUT3 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2023,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_7x: LUT3 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2023,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_m_8x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_M(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_10x: LUT3 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2023,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(10),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_m_11x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(11),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_M(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_m_12x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(12),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_M(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_m_13x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(13),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_M(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_m_14x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(14),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_M(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_m_15x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(15),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_M(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_16x: LUT3 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2023,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(16),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_17x: LUT3 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2023,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_18x: LUT3 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2023,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(18),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_m_21x: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_M(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_22x: LUT3 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2023,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(22),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_23x: LUT3 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2023,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_25x: LUT3 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2023,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(25),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_28x: LUT3 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2023,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(28),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_38x: LUT3 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2023,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(38),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_50x: LUT3 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2023,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(50),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_m_52x: LUT3 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2023,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(52),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_N_2032_i: LUT2 
  generic map(
    INIT => X"E"
  )
  port map (
    I0 => GRLFPC2_0_FPI_START,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(65),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2032_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_112x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(54),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(112),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_506);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_110x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(52),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(110),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_508);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_109x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(109),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_509);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_108x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(50),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(108),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_510);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_107x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(49),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(107),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_511);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_105x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(47),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(105),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_513);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_104x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(46),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(104),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_514);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_103x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(45),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(103),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_515);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_102x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(44),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(102),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_516);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_101x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(43),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(101),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_517);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_93x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(35),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(93),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_525);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_92x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(34),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(92),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_526);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_90x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(32),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(90),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_528);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_88x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(88),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_530);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_82x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(24),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(82),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_536);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_79x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(79),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_539);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_77x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(77),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_541);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_75x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_543);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_74x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(74),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_544);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_73x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(15),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(73),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_545);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_71x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(13),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(71),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_547);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_69x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(11),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(69),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_549);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_68x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(10),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(68),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_550);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_63x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(63),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_555);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_62x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(62),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_556);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_r_sctrl_2_0_0_0x: LUT4_L 
  generic map(
    INIT => X"D8F0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(13),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_2_SN_M1_E_0,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_749);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_86x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(28),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(86),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_532);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_95x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(37),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(95),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_523);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_81x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(81),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_537);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_98x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(98),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_520);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_106x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(48),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(106),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_512);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_87x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(87),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_531);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_85x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(27),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(85),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_533);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_c_pxs_multiplexormulxff_result_0_0_1x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => N_2457,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT0(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_84x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(26),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(84),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_534);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_96x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(38),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(96),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_522);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_78x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(20),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(78),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_540);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_65x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(65),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_553);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_61x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(61),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_557);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_60x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(60),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_558);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_83x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(25),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_535);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_0_91x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(33),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(91),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_527);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_5_sqmuxa: LUT4 
  generic map(
    INIT => X"8000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA_2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(5),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_4_sqmuxa: LUT4 
  generic map(
    INIT => X"40C0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA_2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(5),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_2_sqmuxa_3: LUT4 
  generic map(
    INIT => X"40C0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(5),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_3_sqmuxa_2: LUT4 
  generic map(
    INIT => X"8000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(5),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_55_0: LUT4 
  generic map(
    INIT => X"8CAF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1724,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(57),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_55_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathc_0_1: LUT4 
  generic map(
    INIT => X"AF8C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_0_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_40_0: LUT4 
  generic map(
    INIT => X"AF23"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(56),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_3(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_40_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_54_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(42),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => rfo2_data2(12),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_54_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_35_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(31),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => rfo2_data2(23),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_35_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_41_0: LUT4 
  generic map(
    INIT => X"4C5F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(55),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_41_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_52_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(44),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => rfo2_data2(10),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_52_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_39_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(27),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => rfo2_data2(27),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_39_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_42_0: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(54),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => rfo2_data2(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_42_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_36_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => rfo2_data2(24),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_36_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_19_0: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_19_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_38_0: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(28),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => rfo2_data2(26),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_38_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_46_0: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(50),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => rfo2_data2(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_46_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_44_0: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(52),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => rfo2_data2(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_44_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_43_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(53),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => rfo2_data2(1),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_43_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_14_0: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(22),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(22),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_14_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_13_0: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(23),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(23),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_13_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_12_0: LUT4_L 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(24),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(24),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_12_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_11_0: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(25),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(25),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_11_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_10_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(26),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => rfo2_data2(28),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_10_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_9_0: LUT4 
  generic map(
    INIT => X"4C5F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_9_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_8_0: LUT4 
  generic map(
    INIT => X"4C5F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_8_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_49_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(47),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => rfo2_data2(7),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_49_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_6_0: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(4),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_6_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_5_0: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(5),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_5_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_3_0: LUT3 
  generic map(
    INIT => X"13"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(7),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_3_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_0_0: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(10),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(10),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_0_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_18_0: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(18),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(18),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_18_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_32_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(34),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => rfo2_data2(20),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_32_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_31_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(35),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => rfo2_data2(19),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_31_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_30_0: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(36),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => rfo2_data2(18),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_30_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_29_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(37),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => rfo2_data2(17),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_29_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_28_0: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(38),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => rfo2_data2(16),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_28_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_27_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(39),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => rfo2_data2(15),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_27_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_26_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(40),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => rfo2_data2(14),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_26_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_25_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(41),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => rfo2_data2(13),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_25_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_48_0: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(48),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => rfo2_data2(6),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_48_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_20_0: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(16),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_20_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_17_0: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(19),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1(19),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_17_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un1_xzybus24_s0: LUT2 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un1_xzybus24_s1: LUT2 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_115x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(57),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(115),
    O => N_12496);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_115x: LUT4 
  generic map(
    INIT => X"C0AA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_223,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_ROMXZSL2FROMC,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(118),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => N_12497);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_115x: MUXF5 port map (
      I0 => N_12496,
      I1 => N_12497,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_623);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_113x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(113),
    O => N_12498);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_113x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_223,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_225,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => N_12499);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_113x: MUXF5 port map (
      I0 => N_12498,
      I1 => N_12499,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_625);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_100x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(100),
    O => N_12500);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_100x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(13),
    I1 => GRLFPC2_0_FPO_FRAC(15),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => N_12501);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_100x: MUXF5 port map (
      I0 => N_12500,
      I1 => N_12501,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_638);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_97x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(97),
    O => N_12502);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_97x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(16),
    I1 => GRLFPC2_0_FPO_FRAC(18),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => N_12503);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_97x: MUXF5 port map (
      I0 => N_12502,
      I1 => N_12503,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_641);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_94x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(36),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(94),
    O => N_12504);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_94x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(19),
    I1 => GRLFPC2_0_FPO_FRAC(21),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => N_12505);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_94x: MUXF5 port map (
      I0 => N_12504,
      I1 => N_12505,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_644);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_80x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(22),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(80),
    O => N_12506);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_80x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(33),
    I1 => GRLFPC2_0_FPO_FRAC(35),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => N_12507);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_80x: MUXF5 port map (
      I0 => N_12506,
      I1 => N_12507,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_658);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_76x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(18),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76),
    O => N_12508);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_76x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(37),
    I1 => GRLFPC2_0_FPO_FRAC(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => N_12509);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_76x: MUXF5 port map (
      I0 => N_12508,
      I1 => N_12509,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_662);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_72x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(14),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(72),
    O => N_12510);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_72x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(41),
    I1 => GRLFPC2_0_FPO_FRAC(43),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => N_12511);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_72x: MUXF5 port map (
      I0 => N_12510,
      I1 => N_12511,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_666);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_66x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
    O => N_12512);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_66x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(47),
    I1 => GRLFPC2_0_FPO_FRAC(49),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => N_12513);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_66x: MUXF5 port map (
      I0 => N_12512,
      I1 => N_12513,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_672);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_64x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
    O => N_12514);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_64x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(49),
    I1 => GRLFPC2_0_FPO_FRAC(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => N_12515);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_64x: MUXF5 port map (
      I0 => N_12514,
      I1 => N_12515,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_674);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_59x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(59),
    O => N_12516);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_59x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(54),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_279,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => N_12517);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_59x: MUXF5 port map (
      I0 => N_12516,
      I1 => N_12517,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_679);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_58x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(58),
    O => N_12518);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_58x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_278,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2276,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => N_12519);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_58x: MUXF5 port map (
      I0 => N_12518,
      I1 => N_12519,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_680);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_r_sctrl_3_u_0_am_0x: LUT4 
  generic map(
    INIT => X"CCE4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(13),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_3_SN_I3_I_0,
    O => N_12520);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_r_sctrl_3_u_0_bm_0x: LUT4 
  generic map(
    INIT => X"2772"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2000,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(0),
    I3 => GRLFPC2_0_OP2(63),
    O => N_12521);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_r_sctrl_3_u_0_0x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => N_12520,
    I1 => N_12521,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1529,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_760);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_114x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(56),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(114),
    O => N_12522);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_114x: LUT4 
  generic map(
    INIT => X"C0AA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_224,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_ROMXZSL2FROMC,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(117),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => N_12523);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_114x: MUXF5 port map (
      I0 => N_12522,
      I1 => N_12523,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_624);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_70x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(70),
    O => N_12524);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_70x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(43),
    I1 => GRLFPC2_0_FPO_FRAC(45),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => N_12525);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_70x: MUXF5 port map (
      I0 => N_12524,
      I1 => N_12525,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_668);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_111x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(111),
    O => N_12526);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_111x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(4),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_225,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => N_12527);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_111x: MUXF5 port map (
      I0 => N_12526,
      I1 => N_12527,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_627);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_67x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(9),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(67),
    O => N_12528);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_67x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(46),
    I1 => GRLFPC2_0_FPO_FRAC(48),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => N_12529);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_67x: MUXF5 port map (
      I0 => N_12528,
      I1 => N_12529,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_671);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_99x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(41),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(99),
    O => N_12530);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_99x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(14),
    I1 => GRLFPC2_0_FPO_FRAC(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => N_12531);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_99x: MUXF5 port map (
      I0 => N_12530,
      I1 => N_12531,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_639);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_am_89x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(31),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(89),
    O => N_12532);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_bm_89x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(24),
    I1 => GRLFPC2_0_FPO_FRAC(26),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    O => N_12533);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_3_0_89x: MUXF5 port map (
      I0 => N_12532,
      I1 => N_12533,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_649);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_54_1: LUT3 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_54_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_54_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_52_1: LUT3 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(44),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_52_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_52_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_39_1: LUT3 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(27),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_39_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_39_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_36_1: LUT3 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_36_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_36_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_16_1: LUT4_L 
  generic map(
    INIT => X"0405"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_M(20),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M(20),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(20),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_16_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_15_1: LUT4_L 
  generic map(
    INIT => X"0405"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_M(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M(21),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_15_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_49_1: LUT3 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(47),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_49_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_49_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_4_1: LUT4_L 
  generic map(
    INIT => X"0405"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_M(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M(6),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(6),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_4_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_2_1: LUT4_L 
  generic map(
    INIT => X"0405"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_M(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M(8),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_1_1: LUT4_L 
  generic map(
    INIT => X"0405"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_M(9),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M(9),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(9),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_1_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_1_9: LUT4_L 
  generic map(
    INIT => X"0405"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_M(11),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M(11),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(11),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_22_1: LUT4 
  generic map(
    INIT => X"0405"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_M(14),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M(14),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(14),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_22_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_7_1: LUT4_L 
  generic map(
    INIT => X"0405"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_M(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M(3),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_7_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_29_1: LUT3 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(37),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_29_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_29_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_27_1: LUT3 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_27_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_27_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_26_1: LUT3 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_26_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_26_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_25_1: LUT3 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(41),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_25_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_25_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_24_1: LUT4 
  generic map(
    INIT => X"0405"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_M(12),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M(12),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(12),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_24_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_23_1: LUT4 
  generic map(
    INIT => X"0405"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_M(13),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M(13),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(13),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_23_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_48_1: LUT3 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(48),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_48_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_48_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_21_1: LUT4 
  generic map(
    INIT => X"0405"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_M(15),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M(15),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(15),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_21_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_2_m_54x: LUT4 
  generic map(
    INIT => X"1000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(54),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M(54));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_2_m_53x: LUT4 
  generic map(
    INIT => X"1000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(53),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf0_i_m_55x: LUT3 
  generic map(
    INIT => X"04"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(55),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0_I_M(55));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_notsrres_m_53x: LUT4 
  generic map(
    INIT => X"048C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_1(57),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(53),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(54),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M(53));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_2_m_51x: LUT4 
  generic map(
    INIT => X"1000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(51),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_2_m_48x: LUT4 
  generic map(
    INIT => X"1000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(48),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M(48));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_38x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(38),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(38));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_37x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(37),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(37));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_25x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(25),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(25));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_17x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(17),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(17));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_14x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(14),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf0_m_0x: LUT3 
  generic map(
    INIT => X"40"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0_M(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_0x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf0_m_1x: LUT3 
  generic map(
    INIT => X"40"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0_M(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_2_m_57x: LUT4 
  generic map(
    INIT => X"AC00"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(55),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(57),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_2_m_0_56x: LUT4 
  generic map(
    INIT => X"4000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(56),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M_0(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_2_m_56x: LUT4 
  generic map(
    INIT => X"1000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(56),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M(56));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_2_m_52x: LUT4 
  generic map(
    INIT => X"1000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(52),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M(52));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_2_m_0_51x: LUT4 
  generic map(
    INIT => X"4000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(51),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M_0(51));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_2_m_50x: LUT4 
  generic map(
    INIT => X"1000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(50),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M(50));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_2_m_49x: LUT4 
  generic map(
    INIT => X"1000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(49),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M(49));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_47x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(47),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(47));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_46x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(46),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(46));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_45x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(45),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(45));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_2_m_44x: LUT4 
  generic map(
    INIT => X"AC00"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(42),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(44),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_44x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(44),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_43x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(43),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(43));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_2_m_42x: LUT4 
  generic map(
    INIT => X"AC00"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(40),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_42x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(42),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_41x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(41),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(41));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_40x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(40),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(40));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_39x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(39),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(39));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_36x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(36));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_35x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(35),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(35));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_34x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(34),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(34));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_33x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(33),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(33));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_32x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(32),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(32));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_31x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(31),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(31));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_30x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(30),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(30));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_29x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(29),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(29));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_28x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(28),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(28));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_27x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(27),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(27));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_26x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(26),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(26));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_24x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(24),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(24));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_23x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(23),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(23));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_22x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(22),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(22));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_21x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(21),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(21));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_20x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(20),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_19x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(19),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(19));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_18x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(18),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(18));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_16x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(16),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(16));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_15x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(15),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(15));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_13x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(13),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(13));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_12x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(12),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_11x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(11),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(11));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_10x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(10),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(10));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_9x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(9),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_8x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(8),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_7x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_6x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(6),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_5x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(5),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_4x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_3x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(3),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpuf1_m_2x: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1_M(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_55_2: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(115),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(173),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_55_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathc_1_0: LUT4 
  generic map(
    INIT => X"7030"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_0_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(55),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathc_2_0: LUT4 
  generic map(
    INIT => X"F531"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(60),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(118),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_2_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathc_3: LUT4_L 
  generic map(
    INIT => X"AF23"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(54),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_40_1: LUT4 
  generic map(
    INIT => X"F0B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_40_0,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_40_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_40_2: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(114),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(172),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_40_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_54_3: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(100),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(158),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_54_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_54_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(14),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(43),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_54_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_53_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(101),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(159),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_53_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_51_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(103),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(161),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_51_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_50_2: LUT4 
  generic map(
    INIT => X"F0B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_50_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(11),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_50_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_50_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(104),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(162),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_50_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_50_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(10),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(47),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_50_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_35_2: LUT4 
  generic map(
    INIT => X"F0B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_35_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(26),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_35_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_35_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(89),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(147),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_35_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_35_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(25),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(32),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_35_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_41_1: LUT4 
  generic map(
    INIT => X"F0B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_41_0,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_41_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_41_2: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(113),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(171),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_41_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_41_3: LUT4_L 
  generic map(
    INIT => X"45CF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_224,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2276,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_41_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_52_3: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(102),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(160),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_52_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_52_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(12),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(45),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_52_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_39_2: LUT4 
  generic map(
    INIT => X"F0B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_39_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(30),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_39_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_39_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(85),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(143),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_39_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_39_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(29),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(28),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_39_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_42_2: LUT4 
  generic map(
    INIT => X"0700"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(54),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_42_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_42_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_42_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(112),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(170),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_42_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_42_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_225,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_42_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_37_2: LUT4 
  generic map(
    INIT => X"F0B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_37_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(28),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_37_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_37_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(87),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(145),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_37_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_37_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(27),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(30),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_37_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_36_2: LUT4 
  generic map(
    INIT => X"F0B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_36_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(27),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_36_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_36_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(88),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(146),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_36_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_36_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(26),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(31),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_36_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_19_2: LUT4 
  generic map(
    INIT => X"0700"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_19_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_19_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_19_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(133),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_19_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_19_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(39),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(18),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_19_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_38_2: LUT4 
  generic map(
    INIT => X"0700"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(28),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_38_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_38_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_38_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(86),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(144),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_38_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_38_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(28),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(29),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_38_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_46_2: LUT4 
  generic map(
    INIT => X"0700"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(50),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_46_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_46_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_46_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(108),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(166),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_46_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_46_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_46_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_45_2: LUT4 
  generic map(
    INIT => X"F0B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_45_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(6),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_45_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_45_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(109),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(167),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_45_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_45_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(5),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(52),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_45_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_44_2: LUT4 
  generic map(
    INIT => X"0700"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(52),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_44_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_44_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_44_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(110),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(168),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_44_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_44_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(4),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_44_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_43_2: LUT4 
  generic map(
    INIT => X"F0B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_43_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_43_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_43_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(111),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(169),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_43_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_43_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(54),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_43_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_16_2: LUT4 
  generic map(
    INIT => X"F0B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_16_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(37),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_16_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_16_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(78),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(136),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_16_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_16_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(36),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(21),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_16_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_15_2: LUT4 
  generic map(
    INIT => X"F0B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_15_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_15_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_15_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(79),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(137),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_15_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_15_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(35),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(22),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_15_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_14_2: LUT4 
  generic map(
    INIT => X"0700"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(35),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(22),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_14_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_14_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_14_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(80),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(138),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_14_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_14_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(34),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(23),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_14_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_13_2: LUT4 
  generic map(
    INIT => X"0700"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(34),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(23),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_13_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_13_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_13_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(81),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(139),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_13_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_13_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(33),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(24),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_13_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_12_2: LUT4 
  generic map(
    INIT => X"F0B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_12_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(33),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_12_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_12_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(82),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(140),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_12_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_12_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(32),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(25),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_12_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_11_2: LUT4 
  generic map(
    INIT => X"0700"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(32),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(25),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_11_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_11_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_11_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(141),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_11_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_11_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(31),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(26),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_11_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_10_2: LUT4 
  generic map(
    INIT => X"F0B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_10_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(31),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_10_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_10_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(84),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(142),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_10_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_10_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(27),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_10_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_9_2: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(116),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_9_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_8_2: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(2),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(117),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_8_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_47_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(107),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(165),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_47_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_49_2: LUT4 
  generic map(
    INIT => X"F0B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_49_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(10),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_49_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_49_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(105),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(163),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_49_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_49_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(9),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(48),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_49_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_6_2: LUT4 
  generic map(
    INIT => X"0700"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(62),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(4),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_6_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_6_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_6_3: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(120),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_6_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_34_2: LUT4 
  generic map(
    INIT => X"F0B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_34_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(25),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_34_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_34_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(90),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(148),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_34_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_34_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(24),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(33),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_34_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_33_2: LUT4 
  generic map(
    INIT => X"F0B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_33_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(24),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_33_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_33_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(91),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(149),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_33_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_33_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(34),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_33_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_5_2: LUT4 
  generic map(
    INIT => X"0700"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(63),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(5),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_5_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_5_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_5_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(6),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(121),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_5_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_4_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(7),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(122),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_4_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_3_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(123),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_3_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_2_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(9),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(124),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_2_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_1_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(10),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(125),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_1_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_0_2: LUT4 
  generic map(
    INIT => X"0700"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(47),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(10),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_0_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_0_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_0_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(68),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(126),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_0_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_0_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(46),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(11),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_0_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_2_9: LUT4 
  generic map(
    INIT => X"F0B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(46),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_3_9: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(69),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(127),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_4_9: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(45),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(12),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_22_3: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(72),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(130),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_22_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_22_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(42),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(15),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_22_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_18_2: LUT4 
  generic map(
    INIT => X"0700"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(18),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_18_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_18_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_18_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(134),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_18_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_18_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(38),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(19),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_18_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_7_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(119),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_7_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_32_2: LUT4 
  generic map(
    INIT => X"F0B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_32_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(23),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_32_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_32_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(92),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(150),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_32_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_32_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(22),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(35),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_32_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_31_2: LUT4 
  generic map(
    INIT => X"F0B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_31_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(22),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_31_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_31_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(93),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(151),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_31_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_31_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(36),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_31_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_30_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(94),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(152),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_30_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_30_4: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(20),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(37),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_30_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_29_2: LUT4 
  generic map(
    INIT => X"F0B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_29_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(20),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_29_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_29_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(95),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(153),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_29_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_29_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(19),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(38),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_29_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_28_2: LUT4 
  generic map(
    INIT => X"0700"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(19),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(38),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_28_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_28_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_28_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(96),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(154),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_28_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_28_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(18),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(39),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_28_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_27_2: LUT4 
  generic map(
    INIT => X"F0B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_27_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(18),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_27_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_27_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(97),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(155),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_27_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_27_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(17),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(40),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_27_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_26_2: LUT4 
  generic map(
    INIT => X"F0B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_26_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(17),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_26_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_26_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(98),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(156),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_26_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_26_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(16),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(41),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_26_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_25_2: LUT4 
  generic map(
    INIT => X"F0B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_25_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(16),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_25_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_25_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(99),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(157),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_25_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_25_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(15),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(42),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_25_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_24_3: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(70),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(128),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_24_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_24_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(44),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(13),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_24_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_23_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(71),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(129),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_23_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_23_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(43),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(14),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_23_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_48_3: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(106),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(164),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_48_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_48_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(49),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_48_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_21_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(73),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(131),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_21_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_21_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(41),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(16),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_21_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_20_2: LUT4 
  generic map(
    INIT => X"0700"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(41),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(16),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_20_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_20_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_20_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(74),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(132),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_20_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_20_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(40),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_20_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_17_2: LUT4 
  generic map(
    INIT => X"0700"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(38),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(19),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_17_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_17_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_17_3: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_4_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(77),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(135),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_17_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_17_4: LUT4_L 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(37),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(20),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_17_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_am_112x: LUT4 
  generic map(
    INIT => X"2722"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1752,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I3 => rfo2_data1(0),
    O => N_12534);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_bm_112x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_506,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_566,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12535);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_112x: MUXF5 port map (
      I0 => N_12534,
      I1 => N_12535,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(112));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_am_110x: LUT4 
  generic map(
    INIT => X"2722"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1754,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I3 => rfo2_data1(2),
    O => N_12536);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_bm_110x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_508,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_568,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12537);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_110x: MUXF5 port map (
      I0 => N_12536,
      I1 => N_12537,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(110));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_am_109x: LUT4 
  generic map(
    INIT => X"2722"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1755,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I3 => rfo2_data1(3),
    O => N_12538);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_bm_109x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_509,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_569,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12539);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_109x: MUXF5 port map (
      I0 => N_12538,
      I1 => N_12539,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(109));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_am_108x: LUT4 
  generic map(
    INIT => X"2722"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1756,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I3 => rfo2_data1(4),
    O => N_12540);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_bm_108x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_510,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_570,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12541);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_108x: MUXF5 port map (
      I0 => N_12540,
      I1 => N_12541,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(108));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_am_107x: LUT4 
  generic map(
    INIT => X"2722"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1757,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I3 => rfo2_data1(5),
    O => N_12542);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_bm_107x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_511,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_571,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12543);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_107x: MUXF5 port map (
      I0 => N_12542,
      I1 => N_12543,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(107));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_am_105x: LUT4 
  generic map(
    INIT => X"2722"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1759,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I3 => rfo2_data1(7),
    O => N_12544);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_bm_105x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_513,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_573,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12545);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_105x: MUXF5 port map (
      I0 => N_12544,
      I1 => N_12545,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(105));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_am_104x: LUT4 
  generic map(
    INIT => X"2722"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1760,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I3 => rfo2_data1(8),
    O => N_12546);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_bm_104x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_514,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_574,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12547);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_104x: MUXF5 port map (
      I0 => N_12546,
      I1 => N_12547,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(104));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_am_103x: LUT4 
  generic map(
    INIT => X"2722"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1761,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I3 => rfo2_data1(9),
    O => N_12548);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_bm_103x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_515,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_575,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12549);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_103x: MUXF5 port map (
      I0 => N_12548,
      I1 => N_12549,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(103));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_am_102x: LUT4 
  generic map(
    INIT => X"2722"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1762,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I3 => rfo2_data1(10),
    O => N_12550);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_bm_102x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_516,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_576,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12551);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_102x: MUXF5 port map (
      I0 => N_12550,
      I1 => N_12551,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(102));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_am_101x: LUT4 
  generic map(
    INIT => X"2722"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1763,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I3 => rfo2_data1(11),
    O => N_12552);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_bm_101x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_517,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_577,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12553);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_101x: MUXF5 port map (
      I0 => N_12552,
      I1 => N_12553,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(101));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_100x: MUXF6 port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_459,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_638,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(100));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_97x: MUXF6 port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_462,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_641,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(97));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_94x: MUXF6 port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_465,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_644,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(94));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_am_93x: LUT4 
  generic map(
    INIT => X"2722"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1771,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I3 => rfo2_data1(19),
    O => N_12554);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_bm_93x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_525,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_585,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12555);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_93x: MUXF5 port map (
      I0 => N_12554,
      I1 => N_12555,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(93));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_am_92x: LUT4 
  generic map(
    INIT => X"2722"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1772,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I3 => rfo2_data1(20),
    O => N_12556);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_bm_92x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_526,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_586,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12557);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_92x: MUXF5 port map (
      I0 => N_12556,
      I1 => N_12557,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(92));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_am_90x: LUT4 
  generic map(
    INIT => X"2722"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1774,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I3 => rfo2_data1(22),
    O => N_12558);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_bm_90x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_528,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_588,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12559);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_90x: MUXF5 port map (
      I0 => N_12558,
      I1 => N_12559,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(90));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_am_88x: LUT4 
  generic map(
    INIT => X"2722"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1776,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I3 => rfo2_data1(24),
    O => N_12560);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_bm_88x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_530,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_590,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12561);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_88x: MUXF5 port map (
      I0 => N_12560,
      I1 => N_12561,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(88));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_am_82x: LUT3 
  generic map(
    INIT => X"72"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1782,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(82),
    O => N_12562);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_bm_82x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_536,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_596,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12563);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_82x: MUXF5 port map (
      I0 => N_12562,
      I1 => N_12563,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(82));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_80x: MUXF6 port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_479,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_658,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(80));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_am_79x: LUT3 
  generic map(
    INIT => X"72"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1785,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(79),
    O => N_12564);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_bm_79x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_539,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_599,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12565);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_79x: MUXF5 port map (
      I0 => N_12564,
      I1 => N_12565,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(79));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_am_77x: LUT3 
  generic map(
    INIT => X"72"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1787,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(77),
    O => N_12566);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_bm_77x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_541,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_601,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12567);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_77x: MUXF5 port map (
      I0 => N_12566,
      I1 => N_12567,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(77));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_76x: MUXF6 port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_483,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_662,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(76));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_am_75x: LUT3 
  generic map(
    INIT => X"72"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1789,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(75),
    O => N_12568);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_bm_75x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_543,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_603,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12569);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_75x: MUXF5 port map (
      I0 => N_12568,
      I1 => N_12569,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(75));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_am_74x: LUT3 
  generic map(
    INIT => X"72"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1790,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(74),
    O => N_12570);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_bm_74x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_544,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_604,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12571);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_74x: MUXF5 port map (
      I0 => N_12570,
      I1 => N_12571,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(74));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_am_73x: LUT3 
  generic map(
    INIT => X"72"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1791,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(73),
    O => N_12572);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_bm_73x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_545,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_605,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12573);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_73x: MUXF5 port map (
      I0 => N_12572,
      I1 => N_12573,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(73));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_72x: MUXF6 port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_487,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_666,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(72));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_am_71x: LUT3 
  generic map(
    INIT => X"72"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1793,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(71),
    O => N_12574);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_bm_71x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_547,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_607,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12575);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_71x: MUXF5 port map (
      I0 => N_12574,
      I1 => N_12575,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(71));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_am_69x: LUT3 
  generic map(
    INIT => X"72"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1795,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(69),
    O => N_12576);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_bm_69x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_549,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_609,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12577);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_69x: MUXF5 port map (
      I0 => N_12576,
      I1 => N_12577,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(69));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_am_68x: LUT3 
  generic map(
    INIT => X"72"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1796,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(68),
    O => N_12578);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_bm_68x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_550,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_610,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12579);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_68x: MUXF5 port map (
      I0 => N_12578,
      I1 => N_12579,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(68));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_66x: MUXF6 port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_493,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_672,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(66));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_64x: MUXF6 port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_495,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_674,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(64));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_am_63x: LUT3 
  generic map(
    INIT => X"72"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1801,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(63),
    O => N_12580);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_bm_63x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_555,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_615,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12581);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_63x: MUXF5 port map (
      I0 => N_12580,
      I1 => N_12581,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(63));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_am_62x: LUT3 
  generic map(
    INIT => X"72"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1802,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(62),
    O => N_12582);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_bm_62x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_556,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_616,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12583);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_62x: MUXF5 port map (
      I0 => N_12582,
      I1 => N_12583,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(62));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_am_86x: LUT4 
  generic map(
    INIT => X"2722"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1778,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I3 => rfo2_data1(26),
    O => N_12584);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_bm_86x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_532,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_592,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12585);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_86x: MUXF5 port map (
      I0 => N_12584,
      I1 => N_12585,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(86));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_am_95x: LUT4 
  generic map(
    INIT => X"2722"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1769,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I3 => rfo2_data1(17),
    O => N_12586);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_bm_95x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_523,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_583,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12587);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_95x: MUXF5 port map (
      I0 => N_12586,
      I1 => N_12587,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(95));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_am_81x: LUT3 
  generic map(
    INIT => X"72"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1783,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(81),
    O => N_12588);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_bm_81x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_537,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_597,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12589);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_81x: MUXF5 port map (
      I0 => N_12588,
      I1 => N_12589,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(81));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_am_98x: LUT4 
  generic map(
    INIT => X"2722"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1766,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I3 => rfo2_data1(14),
    O => N_12590);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_bm_98x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_520,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_580,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12591);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_98x: MUXF5 port map (
      I0 => N_12590,
      I1 => N_12591,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(98));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_am_106x: LUT4 
  generic map(
    INIT => X"2722"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1758,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I3 => rfo2_data1(6),
    O => N_12592);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_bm_106x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_512,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_572,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12593);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_106x: MUXF5 port map (
      I0 => N_12592,
      I1 => N_12593,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(106));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_am_87x: LUT4 
  generic map(
    INIT => X"2722"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1777,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I3 => rfo2_data1(25),
    O => N_12594);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_bm_87x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_531,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_591,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12595);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_87x: MUXF5 port map (
      I0 => N_12594,
      I1 => N_12595,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(87));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_am_85x: LUT4 
  generic map(
    INIT => X"2722"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1779,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I3 => rfo2_data1(27),
    O => N_12596);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_bm_85x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_533,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_593,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12597);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_85x: MUXF5 port map (
      I0 => N_12596,
      I1 => N_12597,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(85));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_70x: MUXF6 port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_489,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_668,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(70));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_am_84x: LUT4 
  generic map(
    INIT => X"2722"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1780,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I3 => rfo2_data1(28),
    O => N_12598);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_bm_84x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_534,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_594,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12599);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_84x: MUXF5 port map (
      I0 => N_12598,
      I1 => N_12599,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(84));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_111x: MUXF6 port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_448,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_627,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(111));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_67x: MUXF6 port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_492,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_671,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(67));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_am_96x: LUT4 
  generic map(
    INIT => X"2722"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1768,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I3 => rfo2_data1(16),
    O => N_12600);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_bm_96x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_522,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_582,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12601);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_96x: MUXF5 port map (
      I0 => N_12600,
      I1 => N_12601,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(96));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_99x: MUXF6 port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_460,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_639,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(99));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_89x: MUXF6 port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_470,
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_649,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(89));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_am_78x: LUT3 
  generic map(
    INIT => X"72"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1786,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(78),
    O => N_12602);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_bm_78x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_540,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_600,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12603);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_78x: MUXF5 port map (
      I0 => N_12602,
      I1 => N_12603,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(78));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_am_65x: LUT3 
  generic map(
    INIT => X"72"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1799,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(65),
    O => N_12604);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_bm_65x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_553,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_613,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12605);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_65x: MUXF5 port map (
      I0 => N_12604,
      I1 => N_12605,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(65));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_am_61x: LUT3 
  generic map(
    INIT => X"72"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1803,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(61),
    O => N_12606);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_bm_61x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_557,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_617,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12607);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_61x: MUXF5 port map (
      I0 => N_12606,
      I1 => N_12607,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(61));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_am_60x: LUT4 
  generic map(
    INIT => X"F775"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1812,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_117(52),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_CIN_2,
    O => N_12608);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_bm_60x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_558,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_618,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12609);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_60x: MUXF5 port map (
      I0 => N_12608,
      I1 => N_12609,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_am_83x: LUT3 
  generic map(
    INIT => X"72"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1781,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_19(83),
    O => N_12610);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_bm_83x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_535,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_595,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12611);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_83x: MUXF5 port map (
      I0 => N_12610,
      I1 => N_12611,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(83));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_am_91x: LUT4 
  generic map(
    INIT => X"2722"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1773,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I3 => rfo2_data1(21),
    O => N_12612);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_bm_91x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_527,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_587,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740,
    O => N_12613);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_91x: MUXF5 port map (
      I0 => N_12612,
      I1 => N_12613,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_741,
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(91));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathc_5: LUT3_L 
  generic map(
    INIT => X"70"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(54),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathc_6: LUT4 
  generic map(
    INIT => X"5F13"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(55),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(55),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_40_5: LUT4 
  generic map(
    INIT => X"153F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_40_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_54_5: LUT4_L 
  generic map(
    INIT => X"7000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(15),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_54_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_54_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_54_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_50_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(10),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_50_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_50_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_50_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(11),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(11),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_50_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_35_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(25),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_35_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_35_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_35_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(26),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(26),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_35_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_41_5: LUT3_L 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_41_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2(1),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_41_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_41_6: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_41_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_52_5: LUT4_L 
  generic map(
    INIT => X"7000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(13),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_52_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_52_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_52_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_39_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(29),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_39_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_39_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_39_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(30),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_39_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_42_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_42_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_42_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_42_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(3),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_42_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_37_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(27),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_37_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_37_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_37_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(28),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(28),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_37_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_36_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(26),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_36_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_36_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_36_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(27),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(27),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_36_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_19_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(39),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_19_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_19_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_19_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(40),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(40),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_19_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_38_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(28),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_38_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_38_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_38_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(29),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(29),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_38_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_46_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_46_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_46_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_46_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(7),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_46_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_45_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(5),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_45_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_45_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_45_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(6),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_45_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_44_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(4),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_44_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_44_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_44_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(5),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(5),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_44_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_43_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_43_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_43_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_43_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(4),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(4),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_43_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_16_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(36),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_16_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_16_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_16_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(37),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(37),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_16_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_15_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(35),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_15_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_15_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_15_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(36),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_15_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_14_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(34),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_14_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_14_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_14_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(35),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(35),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_14_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_13_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(33),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_13_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_13_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_13_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(34),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(34),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_13_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_12_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(32),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_12_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_12_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_12_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(33),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(33),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_12_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_11_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(31),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_11_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_11_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_11_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(32),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(32),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_11_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_10_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_10_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_10_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_10_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(31),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(31),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_10_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_9_5: LUT4 
  generic map(
    INIT => X"37BF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(57),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(57),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_9_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_8_5: LUT4 
  generic map(
    INIT => X"37BF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(56),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_8_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_49_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(9),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_49_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_49_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_49_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(10),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(10),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_49_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_6_6: LUT4 
  generic map(
    INIT => X"37BF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(53),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(53),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_6_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_34_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(24),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_34_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_34_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_34_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(25),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(25),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_34_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_33_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_33_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_33_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_33_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(24),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(24),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_33_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_5_6: LUT4 
  generic map(
    INIT => X"37BF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(52),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(52),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_5_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_4_6: LUT4 
  generic map(
    INIT => X"37BF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(51),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(51),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_4_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_3_6: LUT4 
  generic map(
    INIT => X"37BF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(50),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(50),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_3_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_2_6: LUT4 
  generic map(
    INIT => X"37BF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(49),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(49),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_2_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_1_6: LUT4 
  generic map(
    INIT => X"37BF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(48),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(48),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_1_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_0_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(46),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_0_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_0_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_0_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(47),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(47),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_0_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_6_9: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(45),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_7_0: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(46),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(46),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_22_5: LUT4_L 
  generic map(
    INIT => X"7000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(43),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_22_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_22_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_22_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_18_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(38),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_18_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_18_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_18_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(39),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(39),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_18_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_7_6: LUT4 
  generic map(
    INIT => X"37BF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(54),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(54),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_7_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_32_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(22),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_32_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_32_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_32_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(23),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_32_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_31_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_31_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_31_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_31_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(22),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(22),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_31_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_30_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(21),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_30_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_29_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(19),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_29_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_29_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_29_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(20),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(20),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_29_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_28_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(18),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_28_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_28_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_28_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(19),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(19),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_28_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_27_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(17),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_27_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_27_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_27_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(18),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(18),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_27_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_26_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(16),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_26_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_26_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_26_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(17),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(17),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_26_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_25_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(15),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_25_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_25_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_25_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(16),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(16),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_25_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_24_5: LUT4_L 
  generic map(
    INIT => X"7000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(45),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_24_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_24_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_24_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_48_5: LUT4_L 
  generic map(
    INIT => X"7000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(9),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_48_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_48_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_48_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_20_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(40),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_20_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_20_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_20_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(41),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(41),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_20_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_17_6: LUT3_L 
  generic map(
    INIT => X"B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(37),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_17_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_17_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_17_7: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(38),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(38),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_17_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_m_0_am_3x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_76,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1646,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTRESETORUNIMP,
    O => N_12614);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_m_0_bm_3x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => N_2459,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT,
    O => N_12615);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_2_0_6x: MUXF5 port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(6),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_4_2(8),
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_s_2_0_20x: MUXF5 port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(20),
      I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(18),
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
      O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(20));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_31_1: LUT4 
  generic map(
    INIT => X"4F00"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2023,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(35),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_31_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_31_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_32_1: LUT4 
  generic map(
    INIT => X"4F00"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2023,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(34),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_32_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_32_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_10_1: LUT4 
  generic map(
    INIT => X"4F00"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2023,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(26),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_10_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_10_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_12_1: LUT4 
  generic map(
    INIT => X"4F00"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2023,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(24),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_12_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_12_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_43_1: LUT4 
  generic map(
    INIT => X"4F00"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2023,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_43_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_43_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_35_1: LUT4 
  generic map(
    INIT => X"4F00"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2023,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(31),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_35_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_35_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m14_0_am_3x: LUT4 
  generic map(
    INIT => X"0002"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_53_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(9),
    O => N_12164);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_G_57_0: LUT4 
  generic map(
    INIT => X"6696"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(4),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_CIN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(369),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_57_0);
  x_grlfpc2_0_r_mk_rstc: LUT4_L 
  generic map(
    INIT => X"4500"
  )
  port map (
    I0 => GRLFPC2_0_N_710,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1519,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_BUSYMULXFF_UN2_TEMP_3,
    I3 => GRLFPC2_0_R_MK_RSTC_1_0,
    LO => GRLFPC2_0_R_MK_RSTC);
  x_grlfpc2_0_r_mk_ldopc: LUT4_L 
  generic map(
    INIT => X"8000"
  )
  port map (
    I0 => GRLFPC2_0_MOV_7_SQMUXA_3,
    I1 => GRLFPC2_0_R_MK_LDOPC_1,
    I2 => GRLFPC2_0_R_MK_LDOPC_1_0,
    I3 => GRLFPC2_0_R_MK_LDOPC_2,
    LO => GRLFPC2_0_R_MK_LDOPC);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_0_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_0_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_0_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_0_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_0_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_0_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathc: LUT4_L 
  generic map(
    INIT => X"8000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_2_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_5,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_6,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_10_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_10_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_10_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_10_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_10_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_10_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_11_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_11_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_11_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_11_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_11_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_11_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_12_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_12_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_12_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_12_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_12_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_12_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_13_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_13_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_13_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_13_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_13_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_13_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_14_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_14_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_14_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_14_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_14_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_14_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_15_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_15_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_15_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_15_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_15_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_15_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_16_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_16_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_16_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_16_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_16_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_16_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_17_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_17_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_17_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_17_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_17_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_17_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_18_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_18_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_18_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_18_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_18_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_18_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_19_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_19_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_19_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_19_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_19_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_19_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_20_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_20_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_20_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_20_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_20_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_20_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_25_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_25_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_25_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_25_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_25_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_25_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_26_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_26_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_26_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_26_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_26_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_26_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_27_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_27_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_27_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_27_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_27_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_27_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_28_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_28_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_28_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_28_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_28_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_28_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_29_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_29_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_29_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_29_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_29_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_29_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_31_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_31_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_31_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_31_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_31_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_31_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_32_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_32_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_32_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_32_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_32_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_32_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_33_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_33_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_33_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_33_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_33_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_33_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_34_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_34_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_34_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_34_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_34_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_34_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_35_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_35_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_35_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_35_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_35_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_35_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_36_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_36_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_36_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_36_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_36_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_36_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_37_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_37_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_37_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_37_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_37_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_37_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_38_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_38_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_38_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_38_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_38_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_38_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_39_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_39_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_39_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_39_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_39_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_39_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_41_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_41_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_41_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_41_5,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_41_6,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_41_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_42_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_42_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_42_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_42_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_42_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_42_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_43_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_43_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_43_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_43_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_43_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_43_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_44_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_44_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_44_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_44_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_44_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_44_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_45_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_45_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_45_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_45_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_45_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_45_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_46_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_46_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_46_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_46_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_46_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_46_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_49_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_49_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_49_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_49_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_49_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_49_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_50_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_50_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_50_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_50_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_50_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_50_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_N_8703_i: LUT4_L 
  generic map(
    INIT => X"EAC0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW86,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(116),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(118),
    LO => N_8703_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathc_0: LUT3_L 
  generic map(
    INIT => X"20"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_623,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_2_0,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_57_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_57_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(42),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_57_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_58_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_58_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(43),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_58_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_59_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_59_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(44),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_59_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_60_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_60_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(45),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_60_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_61_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_61_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(46),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_61_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_62_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_62_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(47),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_62_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_N_8687_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_63_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(48),
    LO => N_8687_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_N_8702_i: LUT4_L 
  generic map(
    INIT => X"EAC0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW86,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(124),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(126),
    LO => N_8702_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_N_8691_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_65_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(50),
    LO => N_8691_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_N_8701_i: LUT4_L 
  generic map(
    INIT => X"EAC0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW86,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(122),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(124),
    LO => N_8701_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_N_8690_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_67_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(52),
    LO => N_8690_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_N_8700_i: LUT4_L 
  generic map(
    INIT => X"EAC0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW86,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(120),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(122),
    LO => N_8700_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_69_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_69_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(54),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_69_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_70_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_70_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(55),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_70_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_71_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_71_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(56),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_71_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_72_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_72_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(27),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_72_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_N_8689_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_73_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(28),
    LO => N_8689_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_74_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_74_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(29),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_74_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_75_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_75_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(30),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_75_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_76_i: LUT3_L 
  generic map(
    INIT => X"8F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW86,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(142),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_76_0,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_76_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_N_8688_i: LUT4_L 
  generic map(
    INIT => X"8FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW86,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(141),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_77_0,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_77_1,
    LO => N_8688_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_78_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_78_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(33),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_78_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_N_8693_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_79_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(34),
    LO => N_8693_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_80_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_80_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(35),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_80_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_81_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_81_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(36),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_81_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_82_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_82_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(37),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_82_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_83_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_83_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(38),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_83_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_84_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_84_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(39),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_84_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_85_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_85_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(40),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_85_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_86_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_86_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(41),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_86_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_N_8692_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S1_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_87_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(12),
    LO => N_8692_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_88_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_88_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(13),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_88_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_89_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_89_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(14),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_89_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_90_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_90_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(15),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_90_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_91_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_91_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(16),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_91_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_92_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_92_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(17),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_92_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_93_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_93_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(18),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_93_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_94_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_94_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(19),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_94_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_95_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_95_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(20),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_95_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_96_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_96_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(21),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_96_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_97_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_97_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(22),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_97_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_98_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_98_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(23),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_98_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_99_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_99_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(24),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_99_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_N_8699_i: LUT4_L 
  generic map(
    INIT => X"F888"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(25),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2354,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLCREGXZ_XZCREGLOADEN,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(150),
    LO => N_8699_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_101_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_101_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(26),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_101_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_102_i: LUT4_L 
  generic map(
    INIT => X"A820"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2354,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(0),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_102_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_N_8694_i: LUT3_L 
  generic map(
    INIT => X"8F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW86,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(172),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_103_0,
    LO => N_8694_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_104_i: LUT3_L 
  generic map(
    INIT => X"8F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW86,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(171),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_104_0,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_104_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_105_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_105_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(3),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_105_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_106_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_106_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(4),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_106_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_107_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_107_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(5),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_107_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_108_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_108_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(6),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_108_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_109_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_109_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(7),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_109_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_110_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_110_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(8),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_110_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_111_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_111_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(9),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_111_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_112_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_112_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(10),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_112_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_113_i: LUT3_L 
  generic map(
    INIT => X"B3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_113_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(11),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_113_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathc_1: LUT2_L 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_428,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_2_0,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathc_2: LUT4_L 
  generic map(
    INIT => X"C0A0"
  )
  port map (
    I0 => N_2477,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_415,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_2_0,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_N_4,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHC_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_divmultv_0_a2_0x: LUT4_L 
  generic map(
    INIT => X"0002"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(2),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(3),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2297);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_375x: LUT4_L 
  generic map(
    INIT => X"0040"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(3),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_TZ(375),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_I(375));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_115_i: LUT4_L 
  generic map(
    INIT => X"7C3C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(3),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_TZ(375),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_115_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_rndmodeselect_N_1748_i: LUT4_L 
  generic map(
    INIT => X"EFEE"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN1_TEMP,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(2),
    I3 => GRLFPC2_0_R_FSR_RD(1),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1748_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_rndmodeselect_un20_u_rdn_i: LUT4_L 
  generic map(
    INIT => X"FFF4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(21),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(1),
    I3 => GRLFPC2_0_R_FSR_RD(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_RNDMODESELECT_UN20_U_RDN_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_mapmulxff_unimpmap: LUT4_L 
  generic map(
    INIT => X"2103"
  )
  port map (
    I0 => cpi_d_inst(9),
    I1 => cpi_d_inst(13),
    I2 => cpi_d_inst(19),
    I3 => GRLFPC2_0_COMB_FPDECODE_MOV6_2,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW);
  x_grlfpc2_0_comb_v_i_res_1_0_35x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN2_HOLDN,
    I1 => GRLFPC2_0_COMB_V_I_RES_3(35),
    I2 => GRLFPC2_0_OP2(38),
    LO => GRLFPC2_0_COMB_V_I_RES_1(35));
  x_grlfpc2_0_comb_v_i_res_1_0_33x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN2_HOLDN,
    I1 => GRLFPC2_0_COMB_V_I_RES_3(33),
    I2 => GRLFPC2_0_OP2(36),
    LO => GRLFPC2_0_COMB_V_I_RES_1(33));
  x_grlfpc2_0_comb_v_i_res_1_0_32x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN2_HOLDN,
    I1 => GRLFPC2_0_COMB_V_I_RES_3(32),
    I2 => GRLFPC2_0_OP2(35),
    LO => GRLFPC2_0_COMB_V_I_RES_1(32));
  x_grlfpc2_0_r_mk_rst2_i: LUT1_L 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => GRLFPC2_0_R_MK_RST2,
    LO => GRLFPC2_0_R_MK_RST2_I);
  x_grlfpc2_0_comb_v_e_afq_1: LUT3_L 
  generic map(
    INIT => X"10"
  )
  port map (
    I0 => cpi_a_annul,
    I1 => cpi_a_trap,
    I2 => GRLFPC2_0_R_A_AFQ,
    LO => GRLFPC2_0_COMB_V_E_AFQ_1);
  x_grlfpc2_0_comb_v_e_afsr_1: LUT3_L 
  generic map(
    INIT => X"10"
  )
  port map (
    I0 => cpi_a_annul,
    I1 => cpi_a_trap,
    I2 => GRLFPC2_0_R_A_AFSR,
    LO => GRLFPC2_0_COMB_V_E_AFSR_1);
  x_grlfpc2_0_comb_v_e_fpop_1: LUT3_L 
  generic map(
    INIT => X"10"
  )
  port map (
    I0 => cpi_a_annul,
    I1 => cpi_a_trap,
    I2 => GRLFPC2_0_R_A_FPOP,
    LO => GRLFPC2_0_COMB_V_E_FPOP_1);
  x_grlfpc2_0_comb_v_e_ld_1: LUT3_L 
  generic map(
    INIT => X"10"
  )
  port map (
    I0 => cpi_a_annul,
    I1 => cpi_a_trap,
    I2 => GRLFPC2_0_R_A_LD,
    LO => GRLFPC2_0_COMB_V_E_LD_1);
  x_grlfpc2_0_comb_v_m_afq_1: LUT3_L 
  generic map(
    INIT => X"10"
  )
  port map (
    I0 => cpi_e_annul,
    I1 => cpi_e_trap,
    I2 => GRLFPC2_0_R_E_AFQ,
    LO => GRLFPC2_0_COMB_V_M_AFQ_1);
  x_grlfpc2_0_comb_v_m_afsr_1: LUT3_L 
  generic map(
    INIT => X"10"
  )
  port map (
    I0 => cpi_e_annul,
    I1 => cpi_e_trap,
    I2 => GRLFPC2_0_R_E_AFSR,
    LO => GRLFPC2_0_COMB_V_M_AFSR_1);
  x_grlfpc2_0_comb_v_m_fpop_1: LUT3_L 
  generic map(
    INIT => X"10"
  )
  port map (
    I0 => cpi_e_annul,
    I1 => cpi_e_trap,
    I2 => GRLFPC2_0_R_E_FPOP,
    LO => GRLFPC2_0_COMB_V_M_FPOP_1);
  x_grlfpc2_0_comb_v_m_ld_1: LUT3_L 
  generic map(
    INIT => X"10"
  )
  port map (
    I0 => cpi_e_annul,
    I1 => cpi_e_trap,
    I2 => GRLFPC2_0_R_E_LD,
    LO => GRLFPC2_0_COMB_V_M_LD_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_N_1999_i: LUT4_L 
  generic map(
    INIT => X"4044"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(38),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(40),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(13),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1999_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_N_1998_i: LUT4_L 
  generic map(
    INIT => X"4440"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(38),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(40),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(13),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1998_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_Excep_1_4x: LUT4_L 
  generic map(
    INIT => X"00C8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(38),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(40),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_I(41),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1996_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_Excep_1_3x: LUT3_L 
  generic map(
    INIT => X"02"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(38),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(40),
    LO => GRLFPC2_0_FPO_EXC(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_Excep_1_2x: LUT4_L 
  generic map(
    INIT => X"0400"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1990,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(38),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(39),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(40),
    LO => GRLFPC2_0_FPO_EXC(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_Excep_1_1x: LUT4_L 
  generic map(
    INIT => X"0800"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(38),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(39),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(40),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_I(41),
    LO => GRLFPC2_0_FPO_EXC(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_N_1990_i: LUT1_L 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1990,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1990_I);
  x_grlfpc2_0_mov_5_sqmuxa: LUT4_L 
  generic map(
    INIT => X"7000"
  )
  port map (
    I0 => cpi_d_inst(7),
    I1 => cpi_d_inst(8),
    I2 => GRLFPC2_0_COMB_FPDECODE_MOV11,
    I3 => GRLFPC2_0_MOV_5_SQMUXA_2,
    LO => GRLFPC2_0_MOV_5_SQMUXA);
  x_grlfpc2_0_I_245: LUT4_L 
  generic map(
    INIT => X"5044"
  )
  port map (
    I0 => GRLFPC2_0_N_691,
    I1 => GRLFPC2_0_R_I_RDD,
    I2 => GRLFPC2_0_R_X_RDD,
    I3 => GRLFPC2_0_V_I_EXEC_0_SQMUXA,
    LO => GRLFPC2_0_N_692);
  x_grlfpc2_0_comb_v_fsr_nonstd_1_0_0: LUT4_L 
  generic map(
    INIT => X"AC00"
  )
  port map (
    I0 => cpi_dbg_data(22),
    I1 => GRLFPC2_0_COMB_V_FSR_NONSTD_1_M1,
    I2 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
    I3 => rst,
    LO => GRLFPC2_0_COMB_V_FSR_NONSTD_1);
  x_grlfpc2_0_comb_v_fsr_rd_1_0_1x: LUT4_L 
  generic map(
    INIT => X"AC00"
  )
  port map (
    I0 => cpi_dbg_data(31),
    I1 => GRLFPC2_0_COMB_V_FSR_RD_1_M1(1),
    I2 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
    I3 => rst,
    LO => GRLFPC2_0_COMB_V_FSR_RD_1(1));
  x_grlfpc2_0_comb_v_fsr_rd_1_0_0x: LUT4_L 
  generic map(
    INIT => X"AC00"
  )
  port map (
    I0 => cpi_dbg_data(30),
    I1 => GRLFPC2_0_COMB_V_FSR_RD_1_M1(0),
    I2 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
    I3 => rst,
    LO => GRLFPC2_0_COMB_V_FSR_RD_1(0));
  x_grlfpc2_0_comb_v_fsr_tem_1_0_4x: LUT4_L 
  generic map(
    INIT => X"AC00"
  )
  port map (
    I0 => cpi_dbg_data(27),
    I1 => GRLFPC2_0_COMB_V_FSR_TEM_1_M1(4),
    I2 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
    I3 => rst,
    LO => GRLFPC2_0_COMB_V_FSR_TEM_1(4));
  x_grlfpc2_0_comb_v_fsr_tem_1_0_3x: LUT4_L 
  generic map(
    INIT => X"AC00"
  )
  port map (
    I0 => cpi_dbg_data(26),
    I1 => GRLFPC2_0_COMB_V_FSR_TEM_1_M1(3),
    I2 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
    I3 => rst,
    LO => GRLFPC2_0_COMB_V_FSR_TEM_1(3));
  x_grlfpc2_0_comb_v_fsr_tem_1_0_2x: LUT4_L 
  generic map(
    INIT => X"AC00"
  )
  port map (
    I0 => cpi_dbg_data(25),
    I1 => GRLFPC2_0_COMB_V_FSR_TEM_1_M1(2),
    I2 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
    I3 => rst,
    LO => GRLFPC2_0_COMB_V_FSR_TEM_1(2));
  x_grlfpc2_0_comb_v_fsr_tem_1_0_1x: LUT4_L 
  generic map(
    INIT => X"AC00"
  )
  port map (
    I0 => cpi_dbg_data(24),
    I1 => GRLFPC2_0_COMB_V_FSR_TEM_1_M1(1),
    I2 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
    I3 => rst,
    LO => GRLFPC2_0_COMB_V_FSR_TEM_1(1));
  x_grlfpc2_0_comb_v_fsr_tem_1_0_0x: LUT4_L 
  generic map(
    INIT => X"AC00"
  )
  port map (
    I0 => cpi_dbg_data(23),
    I1 => GRLFPC2_0_COMB_V_FSR_TEM_1_M1(0),
    I2 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
    I3 => rst,
    LO => GRLFPC2_0_COMB_V_FSR_TEM_1(0));
  x_grlfpc2_0_comb_v_mk_busy2_2: LUT2_L 
  generic map(
    INIT => X"8"
  )
  port map (
    I0 => GRLFPC2_0_N_710,
    I1 => GRLFPC2_0_R_MK_BUSY,
    LO => GRLFPC2_0_COMB_V_MK_BUSY2_2);
  x_grlfpc2_0_comb_v_mk_busy_2: LUT4_L 
  generic map(
    INIT => X"8A00"
  )
  port map (
    I0 => GRLFPC2_0_N_710,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1519,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_BUSYMULXFF_UN2_TEMP_3,
    I3 => GRLFPC2_0_R_MK_RSTC_1_0,
    LO => GRLFPC2_0_COMB_V_MK_BUSY_2);
  x_grlfpc2_0_comb_N_718_i: LUT3_L 
  generic map(
    INIT => X"BA"
  )
  port map (
    I0 => GRLFPC2_0_N_653,
    I1 => GRLFPC2_0_N_757,
    I2 => GRLFPC2_0_COMB_FPDECODE_AFQ12,
    LO => GRLFPC2_0_N_718_I);
  x_grlfpc2_0_I_237: LUT4_L 
  generic map(
    INIT => X"4000"
  )
  port map (
    I0 => cpi_d_inst(22),
    I1 => cpi_d_inst(31),
    I2 => GRLFPC2_0_I_237_2,
    I3 => GRLFPC2_0_N_703_1,
    LO => GRLFPC2_0_N_703);
  x_grlfpc2_0_N_657_i: LUT4_L 
  generic map(
    INIT => X"EFAA"
  )
  port map (
    I0 => GRLFPC2_0_N_653,
    I1 => GRLFPC2_0_N_654,
    I2 => GRLFPC2_0_N_757,
    I3 => GRLFPC2_0_COMB_FPDECODE_AFQ12,
    LO => GRLFPC2_0_N_657_I);
  x_grlfpc2_0_v_fsr_N_721_i: LUT4_L 
  generic map(
    INIT => X"DC00"
  )
  port map (
    I0 => GRLFPC2_0_N_755,
    I1 => GRLFPC2_0_COMB_V_I_V6,
    I2 => GRLFPC2_0_R_FSR_FTT(0),
    I3 => rst,
    LO => GRLFPC2_0_N_721_I);
  x_grlfpc2_0_v_fsr_N_720_i: LUT4_L 
  generic map(
    INIT => X"F040"
  )
  port map (
    I0 => GRLFPC2_0_N_755,
    I1 => GRLFPC2_0_R_FSR_FTT(2),
    I2 => GRLFPC2_0_V_FSR_FTT_1_SQMUXA_2_1,
    I3 => GRLFPC2_0_V_FSR_FTT_1_SQMUXA_2_2,
    LO => GRLFPC2_0_N_720_I);
  x_grlfpc2_0_I_190: LUT4_L 
  generic map(
    INIT => X"8C04"
  )
  port map (
    I0 => cpi_d_inst(23),
    I1 => cpi_d_inst(31),
    I2 => GRLFPC2_0_N_635,
    I3 => GRLFPC2_0_N_636,
    LO => GRLFPC2_0_N_637);
  x_grlfpc2_0_I_173: LUT4_L 
  generic map(
    INIT => X"BF00"
  )
  port map (
    I0 => GRLFPC2_0_N_653,
    I1 => GRLFPC2_0_N_654,
    I2 => GRLFPC2_0_N_757,
    I3 => GRLFPC2_0_COMB_FPDECODE_AFQ12,
    LO => GRLFPC2_0_N_615);
  x_grlfpc2_0_comb_v_state_1_iv_1x: LUT4_L 
  generic map(
    INIT => X"F800"
  )
  port map (
    I0 => cpi_exack,
    I1 => CPO_EXC_INT_2,
    I2 => GRLFPC2_0_COMB_V_STATE_7(1),
    I3 => GRLFPC2_0_V_STATE_1_SQMUXA,
    LO => GRLFPC2_0_COMB_V_STATE_1(1));
  x_grlfpc2_0_comb_v_state_1_0x: LUT4_L 
  generic map(
    INIT => X"7000"
  )
  port map (
    I0 => cpi_exack,
    I1 => CPO_EXC_INT_2,
    I2 => GRLFPC2_0_COMB_V_STATE_7(0),
    I3 => GRLFPC2_0_V_STATE_1_SQMUXA,
    LO => GRLFPC2_0_COMB_V_STATE_1(0));
  x_grlfpc2_0_comb_v_fsr_fcc_1_0_1x: LUT3_L 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(11),
    I1 => GRLFPC2_0_COMB_V_FSR_FCC_1_M1(1),
    I2 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
    LO => GRLFPC2_0_COMB_V_FSR_FCC_1(1));
  x_grlfpc2_0_comb_v_fsr_fcc_1_0_0x: LUT3_L 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => cpi_dbg_data(10),
    I1 => GRLFPC2_0_COMB_V_FSR_FCC_1_M1(0),
    I2 => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1,
    LO => GRLFPC2_0_COMB_V_FSR_FCC_1(0));
  x_grlfpc2_0_I_162: LUT4_L 
  generic map(
    INIT => X"0008"
  )
  port map (
    I0 => GRLFPC2_0_I_162_1,
    I1 => GRLFPC2_0_N_789,
    I2 => GRLFPC2_0_COMB_CCWR4,
    I3 => GRLFPC2_0_COMB_WRRES4,
    LO => GRLFPC2_0_N_602);
  x_grlfpc2_0_comb_v_fsr_N_728_i: LUT4_L 
  generic map(
    INIT => X"FD55"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_1(4),
    I1 => GRLFPC2_0_R_FSR_AEXC(4),
    I2 => GRLFPC2_0_R_I_EXC(4),
    I3 => GRLFPC2_0_V_FSR_CEXC_0_SQMUXA,
    LO => GRLFPC2_0_N_728_I);
  x_grlfpc2_0_comb_v_fsr_N_729_i: LUT4_L 
  generic map(
    INIT => X"FD55"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_1(3),
    I1 => GRLFPC2_0_R_FSR_AEXC(3),
    I2 => GRLFPC2_0_R_I_EXC(3),
    I3 => GRLFPC2_0_V_FSR_CEXC_0_SQMUXA,
    LO => GRLFPC2_0_N_729_I);
  x_grlfpc2_0_comb_v_fsr_N_730_i: LUT4_L 
  generic map(
    INIT => X"FD55"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_1(2),
    I1 => GRLFPC2_0_R_FSR_AEXC(2),
    I2 => GRLFPC2_0_R_I_EXC(2),
    I3 => GRLFPC2_0_V_FSR_CEXC_0_SQMUXA,
    LO => GRLFPC2_0_N_730_I);
  x_grlfpc2_0_comb_v_fsr_N_731_i: LUT4_L 
  generic map(
    INIT => X"FD55"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_1(1),
    I1 => GRLFPC2_0_R_FSR_AEXC(1),
    I2 => GRLFPC2_0_R_I_EXC(1),
    I3 => GRLFPC2_0_V_FSR_CEXC_0_SQMUXA,
    LO => GRLFPC2_0_N_731_I);
  x_grlfpc2_0_comb_v_fsr_N_732_i: LUT4_L 
  generic map(
    INIT => X"FD55"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_FSR_AEXC_1_IV_1(0),
    I1 => GRLFPC2_0_R_FSR_AEXC(0),
    I2 => GRLFPC2_0_R_I_EXC(0),
    I3 => GRLFPC2_0_V_FSR_CEXC_0_SQMUXA,
    LO => GRLFPC2_0_N_732_I);
  x_grlfpc2_0_comb_v_a_afq_1: LUT3_L 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_AFQ_3_SQMUXA,
    I1 => GRLFPC2_0_R_MK_LDOPC_1,
    I2 => GRLFPC2_0_R_MK_LDOPC_2,
    LO => GRLFPC2_0_COMB_V_A_AFQ_1);
  x_grlfpc2_0_comb_v_a_ld_1: LUT3_L 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_COMB_SEQERR_UN13_OP,
    I1 => GRLFPC2_0_R_MK_LDOPC_1,
    I2 => GRLFPC2_0_R_MK_LDOPC_2,
    LO => GRLFPC2_0_COMB_V_A_LD_1);
  x_grlfpc2_0_comb_v_a_st_1: LUT3_L 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_COMB_FPDECODE_ST,
    I1 => GRLFPC2_0_R_MK_LDOPC_1,
    I2 => GRLFPC2_0_R_MK_LDOPC_2,
    LO => GRLFPC2_0_COMB_V_A_ST_1);
  x_grlfpc2_0_comb_v_i_v_1_f0: LUT4_L 
  generic map(
    INIT => X"50D0"
  )
  port map (
    I0 => GRLFPC2_0_N_762,
    I1 => GRLFPC2_0_R_I_V,
    I2 => GRLFPC2_0_V_I_EXEC26,
    I3 => holdn,
    LO => GRLFPC2_0_COMB_V_I_V_1);
  x_grlfpc2_0_comb_v_a_afsr_1_0: LUT4_L 
  generic map(
    INIT => X"8000"
  )
  port map (
    I0 => GRLFPC2_0_COMB_FPDECODE_AFQ13,
    I1 => GRLFPC2_0_COMB_V_A_AFSR_1_0_1,
    I2 => GRLFPC2_0_R_MK_LDOPC_1,
    I3 => GRLFPC2_0_R_MK_LDOPC_2,
    LO => GRLFPC2_0_COMB_V_A_AFSR_1);
  x_grlfpc2_0_comb_v_a_seqerr_1: LUT3_L 
  generic map(
    INIT => X"40"
  )
  port map (
    I0 => GRLFPC2_0_N_736,
    I1 => GRLFPC2_0_R_MK_LDOPC_1,
    I2 => GRLFPC2_0_R_MK_LDOPC_2,
    LO => GRLFPC2_0_COMB_V_A_SEQERR_1);
  x_grlfpc2_0_comb_rdd_1_0: LUT4_L 
  generic map(
    INIT => X"40CC"
  )
  port map (
    I0 => cpi_d_inst(30),
    I1 => GRLFPC2_0_COMB_RDD_1_0_0,
    I2 => GRLFPC2_0_MOV_2_SQMUXA,
    I3 => GRLFPC2_0_UN1_AFQ7_I_A2_2,
    LO => GRLFPC2_0_COMB_RDD_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_un61_pctrl_new_i: LUT3_L 
  generic map(
    INIT => X"FB"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(61),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP_1,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_UN61_PCTRL_NEW_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_pctrl_new_18_74x: LUT2_L 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(62),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_PCTRL_NEW_18(74));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_startshft_un3_notresetorunimp_i: LUT1_L 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTRESETORUNIMP,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN3_NOTRESETORUNIMP_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_N_1519_i: LUT4_L 
  generic map(
    INIT => X"CFAF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_361,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_372,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_0,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(49),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1519_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_un72_pctrl_new_i: LUT4_L 
  generic map(
    INIT => X"EEAE"
  )
  port map (
    I0 => GRLFPC2_0_FPI_START,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_TEMP_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN1_MIFROMINST_0,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WAITMULXFF_NOTSAMPLEDWAIT,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_UN72_PCTRL_NEW_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_startshft_un2_notdecodedunimp_i: LUT1_L 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN2_NOTDECODEDUNIMP,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN2_NOTDECODEDUNIMP_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_N_1723_i: LUT3_L 
  generic map(
    INIT => X"EF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_STARTSHFT_UN2_NOTDECODEDUNIMP,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(64),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(68),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1723_I);
  x_grlfpc2_0_fpi_N_774_i: LUT2_L 
  generic map(
    INIT => X"7"
  )
  port map (
    I0 => GRLFPC2_0_N_782,
    I1 => rst,
    LO => GRLFPC2_0_N_774_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_resvec_0_0x: LUT3_L 
  generic map(
    INIT => X"A3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(4),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_RESVEC(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_i_42x: LUT1_L 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(42),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_I(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_r_sctrl_1_i_0x: LUT3_L 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(5),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_TEMP,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_SCTRL_1_I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_r_sctrl_2_u_0_0x: LUT3_L 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_749,
    I2 => GRLFPC2_0_OP1(63),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_752);
  x_I_761: LUT1_L 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => cpi_d_inst(6),
    LO => CPI_D_INST_I(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_N_1741_i: LUT4_L 
  generic map(
    INIT => X"BAEA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN1_U_SNNOTDB,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN4_TOGGLESIG,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_UN12_U_SNNOTDB_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1741_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_N_1728_i: LUT4_L 
  generic map(
    INIT => X"2013"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_760,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1741,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8(8),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8(9),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1728_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_sctrl_new_16_6x: LUT3_L 
  generic map(
    INIT => X"01"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1741,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8(9),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_16(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_un109_sctrl_new: LUT2_L 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8(9),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SCTRL_NEW_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_sctrl_new_14_4x: LUT4_L 
  generic map(
    INIT => X"2010"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_760,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1741,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8(8),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8(9),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_14(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_sctrl_new_13_3x: LUT3_L 
  generic map(
    INIT => X"84"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_760,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_8(9),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_13(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_sctrl_new_4_2x: LUT3_L 
  generic map(
    INIT => X"40"
  )
  port map (
    I0 => cpi_d_inst(7),
    I1 => cpi_d_inst(9),
    I2 => GRLFPC2_0_COMB_FPDECODE_MOV6_2,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_4(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_sctrl_new_5_1x: LUT3_L 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => cpi_d_inst(7),
    I1 => cpi_d_inst(9),
    I2 => GRLFPC2_0_COMB_FPDECODE_MOV6_2,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SCTRL_NEW_5(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_sxc_N_1997_i: LUT4_L 
  generic map(
    INIT => X"F200"
  )
  port map (
    I0 => cpi_d_inst(7),
    I1 => cpi_d_inst(8),
    I2 => cpi_d_inst(9),
    I3 => GRLFPC2_0_COMB_FPDECODE_MOV6_2,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1997_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_mixoin_3_i_0x: LUT4_L 
  generic map(
    INIT => X"15D5"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1743,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN42_NOTPROP,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN49_NOTPROP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_2(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_3_I(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1766_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1850,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_155(14),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_14_TRFWWBASICCELL_CIN,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1766_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1765_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1851,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_156(13),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_13_TRFWWBASICCELL_CIN_1,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1765_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1764_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1852,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_157(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_12_TRFWWBASICCELL_CIN,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1764_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1763_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1853,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_158(11),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_11_TRFWWBASICCELL_CIN_2,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1763_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1762_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1854,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_159(10),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_10_TRFWWBASICCELL_CIN_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1762_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1761_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1855,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_160(9),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_9_TRFWWBASICCELL_CIN_2,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1761_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1760_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1856,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_161(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_8_TRFWWBASICCELL_CIN,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1760_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1759_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1857,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_162(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_7_TRFWWBASICCELL_CIN_2,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1759_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1758_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1858,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_163(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_6_TRFWWBASICCELL_CIN,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1758_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1757_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1859,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_164(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_5_TRFWWBASICCELL_CIN,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1757_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1756_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1860,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_165(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_4_TRFWWBASICCELL_CIN,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1756_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1755_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1861,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_166(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_3_TRFWWBASICCELL_CIN_2,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1755_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1754_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1862,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_167(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_2_TRFWWBASICCELL_CIN_2,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1754_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1753_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1863,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_168(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_1_TRFWWBASICCELL_CIN_1,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1753_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1752_i: LUT4_L 
  generic map(
    INIT => X"D540"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1865,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_TEMP2_3,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1752_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1781_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1835,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_140(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_29_TRFWWBASICCELL_CIN_1,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1781_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1780_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1836,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_141(28),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_28_TRFWWBASICCELL_CIN_2,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1780_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1779_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1837,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_142(27),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_27_TRFWWBASICCELL_CIN_2,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1779_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1778_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1838,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_143(26),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_26_TRFWWBASICCELL_CIN_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1778_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1777_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1839,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_144(25),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_25_TRFWWBASICCELL_CIN,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1777_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1776_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1840,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_145(24),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_24_TRFWWBASICCELL_CIN_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1776_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1775_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1841,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_146(23),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_23_TRFWWBASICCELL_CIN_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1775_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1774_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1842,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_147(22),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_22_TRFWWBASICCELL_CIN_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1774_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1773_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1843,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_148(21),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_21_TRFWWBASICCELL_CIN_2,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1773_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1772_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1844,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_149(20),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_20_TRFWWBASICCELL_CIN_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1772_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1771_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1845,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_150(19),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_19_TRFWWBASICCELL_CIN_2,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1771_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1770_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1846,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_151(18),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_18_TRFWWBASICCELL_CIN,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1770_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1769_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1847,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_152(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_17_TRFWWBASICCELL_CIN_2,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1769_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1768_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1848,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_153(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_16_TRFWWBASICCELL_CIN_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1768_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1767_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1849,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_154(15),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_15_TRFWWBASICCELL_CIN_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1767_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1796_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1820,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_125(44),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_44_TRFWWBASICCELL_CIN_1,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1796_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1795_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1821,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_126(43),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_43_TRFWWBASICCELL_CIN_2,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1795_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1794_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1822,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_127(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_42_TRFWWBASICCELL_CIN_2,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1794_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1793_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1823,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_128(41),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_41_TRFWWBASICCELL_CIN_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1793_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1792_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1824,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_129(40),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_40_TRFWWBASICCELL_CIN,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1792_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1791_i: LUT4_L 
  generic map(
    INIT => X"D450"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1825,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_130(39),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_39_TRFWWBASICCELL_TEMP2_2,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1791_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1790_i: LUT4_L 
  generic map(
    INIT => X"D450"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1826,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_131(38),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_38_TRFWWBASICCELL_TEMP2_2,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1790_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1789_i: LUT4_L 
  generic map(
    INIT => X"D450"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1827,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_132(37),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_37_TRFWWBASICCELL_TEMP2_1,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1789_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1788_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1828,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_133(36),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_36_TRFWWBASICCELL_CIN_2,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1788_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1787_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1829,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_134(35),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_35_TRFWWBASICCELL_CIN_1,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1787_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1786_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1830,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_135(34),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_34_TRFWWBASICCELL_CIN_1,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1786_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1785_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1831,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_136(33),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_33_TRFWWBASICCELL_CIN_1,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1785_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1784_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1832,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_137(32),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_32_TRFWWBASICCELL_CIN_2,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1784_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1783_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1833,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_138(31),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_31_TRFWWBASICCELL_CIN_1,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1783_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1782_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1834,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_139(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_30_TRFWWBASICCELL_CIN_1,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1782_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1724_i: LUT4_L 
  generic map(
    INIT => X"FDDD"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_5(57),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN28_STKOUT,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN42_NOTPROP,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_2(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1724_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1751_i: LUT4_L 
  generic map(
    INIT => X"4DD4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1810,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_CIN_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_CIN_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_114_1(56),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1751_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1806_i: LUT4_L 
  generic map(
    INIT => X"4DD4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1810,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_54_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_CIN_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_114_1(56),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1806_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1805_i: LUT4_L 
  generic map(
    INIT => X"4DD4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1811,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_53_TRFWWBASICCELL_CIN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_55_TRFWWBASICCELL_CIN,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_114_1(56),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1805_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_23_i_i_60x: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1812,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_117(52),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_52_TRFWWBASICCELL_CIN_2,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23_I_I(60));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1803_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1813,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_1(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_51_TRFWWBASICCELL_CIN_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1803_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1802_i: LUT4_L 
  generic map(
    INIT => X"71D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1814,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2119,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_50_TRFWWBASICCELL_CIN_2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_SI_114_1_1_0(56),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1802_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1801_i: LUT4_L 
  generic map(
    INIT => X"D741"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1815,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1874,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_120_1(49),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_49_TRFWWBASICCELL_CIN_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1801_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1800_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1816,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_121(48),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_48_TRFWWBASICCELL_CIN_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1800_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1799_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1817,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_122(47),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_47_TRFWWBASICCELL_CIN_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1799_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1798_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1818,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_123(46),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_46_TRFWWBASICCELL_CIN_1,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1798_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_N_1797_i: LUT3_L 
  generic map(
    INIT => X"D4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1819,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_56_SI_124(45),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_45_TRFWWBASICCELL_CIN_1,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1797_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_252x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_382,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_422,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(252));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_253x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_381,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_421,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(253));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_254x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_380,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_420,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(254));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_255x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_379,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_419,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(255));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_256x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_378,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_418,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(256));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_257x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_377,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_417,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(257));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_49_258x: LUT3_L 
  generic map(
    INIT => X"6A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_49_1(258),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_mlogd_UN79_ZERO,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_TRFWWBASICCELL_TEMP2_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_49(258));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_237x: LUT3_L 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_770,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_809,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_815,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(237));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_238x: LUT3_L 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_769,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_808,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_815,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(238));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_239x: LUT3_L 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_768,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_807,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_815,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(239));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_240x: LUT3_L 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_767,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_806,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_815,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(240));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_241x: LUT3_L 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_766,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_805,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_815,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(241));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_242x: LUT3_L 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_765,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_804,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_815,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(242));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_243x: LUT3_L 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_764,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_803,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_815,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(243));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_244x: LUT3_L 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_763,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_802,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_815,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(244));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_247x: LUT4_L 
  generic map(
    INIT => X"8D88"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_427,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I3 => GRLFPC2_0_OP1(62),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(247));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_248x: LUT4_L 
  generic map(
    INIT => X"8D88"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_426,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I3 => GRLFPC2_0_OP1(61),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(248));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_249x: LUT4_L 
  generic map(
    INIT => X"8D88"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_425,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_SCTRL(11),
    I3 => GRLFPC2_0_OP1(60),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(249));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_250x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_384,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_424,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(250));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_251x: LUT3_L 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_383,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_423,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(251));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_113x: LUT4_L 
  generic map(
    INIT => X"A088"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_625,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(113),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(113));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_4_114x: LUT4_L 
  generic map(
    INIT => X"08A8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_624,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_3(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(114));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_58x: LUT4_L 
  generic map(
    INIT => X"0A88"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_680,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1806,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(58));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_1_59x: LUT4_L 
  generic map(
    INIT => X"0A88"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_679,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1805,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(59));
  x_grlfpc2_0_comb_v_fsr_N_727_i_1: LUT4 
  generic map(
    INIT => X"153F"
  )
  port map (
    I0 => cpi_lddata(0),
    I1 => GRLFPC2_0_R_I_EXC(0),
    I2 => GRLFPC2_0_V_FSR_CEXC_0_SQMUXA,
    I3 => GRLFPC2_0_V_FSR_CEXC_2_SQMUXA,
    O => GRLFPC2_0_COMB_V_FSR_N_727_I_1);
  x_grlfpc2_0_comb_v_fsr_N_726_i_1: LUT4 
  generic map(
    INIT => X"153F"
  )
  port map (
    I0 => cpi_lddata(1),
    I1 => GRLFPC2_0_R_I_EXC(1),
    I2 => GRLFPC2_0_V_FSR_CEXC_0_SQMUXA,
    I3 => GRLFPC2_0_V_FSR_CEXC_2_SQMUXA,
    O => GRLFPC2_0_COMB_V_FSR_N_726_I_1);
  x_grlfpc2_0_comb_v_fsr_N_725_i_1: LUT4 
  generic map(
    INIT => X"153F"
  )
  port map (
    I0 => cpi_lddata(2),
    I1 => GRLFPC2_0_R_I_EXC(2),
    I2 => GRLFPC2_0_V_FSR_CEXC_0_SQMUXA,
    I3 => GRLFPC2_0_V_FSR_CEXC_2_SQMUXA,
    O => GRLFPC2_0_COMB_V_FSR_N_725_I_1);
  x_grlfpc2_0_comb_v_fsr_N_724_i_1: LUT4 
  generic map(
    INIT => X"153F"
  )
  port map (
    I0 => cpi_lddata(3),
    I1 => GRLFPC2_0_R_I_EXC(3),
    I2 => GRLFPC2_0_V_FSR_CEXC_0_SQMUXA,
    I3 => GRLFPC2_0_V_FSR_CEXC_2_SQMUXA,
    O => GRLFPC2_0_COMB_V_FSR_N_724_I_1);
  x_grlfpc2_0_comb_v_fsr_N_723_i_1: LUT4 
  generic map(
    INIT => X"153F"
  )
  port map (
    I0 => cpi_lddata(4),
    I1 => GRLFPC2_0_R_I_EXC(4),
    I2 => GRLFPC2_0_V_FSR_CEXC_0_SQMUXA,
    I3 => GRLFPC2_0_V_FSR_CEXC_2_SQMUXA,
    O => GRLFPC2_0_COMB_V_FSR_N_723_I_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_40_i_1: LUT4 
  generic map(
    INIT => X"0777"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_223,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_40_I_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_9_6_1: LUT4 
  generic map(
    INIT => X"135F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_279,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(58),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_9_6_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_25_0_0_1: LUT4 
  generic map(
    INIT => X"03F5"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(51),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(52),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_25_0_0_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_33_1_1: LUT4_L 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(33),
    I3 => rfo2_data2(21),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_33_1_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_33_1: LUT3 
  generic map(
    INIT => X"70"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(33),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_33_1_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_33_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_34_1_1: LUT4_L 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(32),
    I3 => rfo2_data2(22),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_34_1_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_34_1: LUT3 
  generic map(
    INIT => X"70"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(32),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_34_1_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_34_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_47_1_1: LUT4_L 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(49),
    I3 => rfo2_data2(5),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_47_1_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_47_1: LUT3 
  generic map(
    INIT => X"70"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(49),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_47_1_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_47_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_45_1_1: LUT4_L 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
    I3 => rfo2_data2(3),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_45_1_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_45_1: LUT3 
  generic map(
    INIT => X"70"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(51),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_45_1_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_45_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_37_1_1: LUT4_L 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(29),
    I3 => rfo2_data2(25),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_37_1_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_37_1: LUT3 
  generic map(
    INIT => X"70"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(29),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_37_1_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_37_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_50_1_1: LUT4_L 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(46),
    I3 => rfo2_data2(8),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_50_1_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpathsr_50_1: LUT3 
  generic map(
    INIT => X"70"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(46),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_50_1_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_50_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_iv_i_141_223_1: LUT3 
  generic map(
    INIT => X"15"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(374),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(375),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(376),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_IV_I_141_223_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_iv_i_141_223: LUT4 
  generic map(
    INIT => X"02A0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2371,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(375),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(377),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_IV_I_141_223_1,
    O => N_2376);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_35_1: LUT4 
  generic map(
    INIT => X"65A5"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(31),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS24,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_IV_0(31),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(25),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_35_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzZero_1_35: LUT4 
  generic map(
    INIT => X"8008"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN22_XZXBUS_5_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_19,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_35_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1_35);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_notprop_1_1: LUT4 
  generic map(
    INIT => X"7717"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_TRFWWRRAY_REMWmul61_0_TRFWWBASICCELL_CIN_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(370),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_NOTPROP_1_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_mullsblogic_stckypair_notprop_1: LUT4 
  generic map(
    INIT => X"2184"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_G_57_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_SALSBS(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_NOTPROP_1_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_TEMP_1(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1869);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_1_1_57x: LUT4_L 
  generic map(
    INIT => X"6801"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN9_NOTPROP,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_1_1(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_dpath_new_8_1_57x: LUT3 
  generic map(
    INIT => X"A2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_1_1(57),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(315),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8_1(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_mixoin_0_1_0x: LUT3_L 
  generic map(
    INIT => X"17"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(1),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_0_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_mixoin_0_0x: LUT3 
  generic map(
    INIT => X"71"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_SUMIN_4(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_CTRLXERSHFT_MIXOIN_3(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_0_1(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_reexcovuv_un30_locov_1: LUT4 
  generic map(
    INIT => X"017F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_EXP(8),
    I1 => GRLFPC2_0_FPO_EXP(9),
    I2 => GRLFPC2_0_FPO_EXP(10),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN30_LOCOV_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_entryshft_un1_s_14_1: LUT4_L 
  generic map(
    INIT => X"0A30"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_ENTRYSHFT_S_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(80),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(83),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(84),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN1_S_14_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_entryshft_un1_s_14: LUT4_L 
  generic map(
    INIT => X"F531"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN1_S_14_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN9_S_11_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(79),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(81),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_ENTRYSHFT_UN1_S_14);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_reexcovuv_un20_locov_5_1: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_FPO_EXP(1),
    I1 => GRLFPC2_0_FPO_EXP(2),
    I2 => GRLFPC2_0_FPO_EXP(3),
    I3 => GRLFPC2_0_FPO_EXP(4),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN20_LOCOV_5_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_reexcovuv_un20_locov_5: LUT4 
  generic map(
    INIT => X"0080"
  )
  port map (
    I0 => GRLFPC2_0_FPO_EXP(5),
    I1 => GRLFPC2_0_FPO_EXP(6),
    I2 => GRLFPC2_0_FPO_EXP(7),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN20_LOCOV_5_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN20_LOCOV_5);
  x_g2_2: LUT3 
  generic map(
    INIT => X"DF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(47),
    I1 => GRLFPC2_0_R_MK_RST2,
    I2 => rst,
    O => G2_2);
  x_g0_4: LUT4_L 
  generic map(
    INIT => X"0CAC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPYBUS_2(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(237),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    LO => N_12635);
  x_g0_5: LUT4_L 
  generic map(
    INIT => X"0CAC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPYBUS_2(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(236),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
    LO => N_12636);
  x_g2_4: LUT4 
  generic map(
    INIT => X"FFFE"
  )
  port map (
    I0 => G2_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE(12),
    I2 => GRLFPC2_0_R_MK_LDOP,
    I3 => GRLFPC2_0_R_MK_RST,
    O => G2_4);
  x_g0_0_x2: LUT4 
  generic map(
    INIT => X"6C93"
  )
  port map (
    I0 => N_12635,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => N_12633);
  x_g0_0_x2_0: LUT4 
  generic map(
    INIT => X"6C93"
  )
  port map (
    I0 => N_12636,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => N_12634);
  x_g4_2: LUT4 
  generic map(
    INIT => X"0100"
  )
  port map (
    I0 => N_12633,
    I1 => N_12634,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_9,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_NE_4,
    O => G4_2);
  x_g4_5: LUT4 
  generic map(
    INIT => X"0200"
  )
  port map (
    I0 => G4_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_NE_10,
    O => G4_5);
  x_grlfpc2_0_r_x_rdd_0_0_I_1: SRL16E port map (
      Q => GRLFPC2_0_R_X_RDD_0_0_TMP_D_ARRAY_0(0),
      A0 => NN_1,
      A1 => NN_2,
      A2 => NN_1,
      A3 => NN_1,
      D => GRLFPC2_0_COMB_RDD_1,
      CLK => clk,
      CE => holdn);
  x_grlfpc2_0_r_x_seqerr_0_0_I_1: SRL16E port map (
      Q => GRLFPC2_0_R_X_SEQERR_0_0_N_6,
      A0 => NN_1,
      A1 => NN_2,
      A2 => NN_1,
      A3 => NN_1,
      D => GRLFPC2_0_COMB_V_A_SEQERR_1,
      CLK => clk,
      CE => holdn);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_fast_376x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_FAST(376),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2297,
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2298);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_fast_10x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_FAST,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1741_I,
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_10_rep1: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP1,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1741_I,
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_sctrl_10_rep2: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_REP2,
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1741_I,
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_sqmuxa_1_L1_0: LUT2 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(7),
    O => N_12791);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_8_sqmuxa_1: LUT4 
  generic map(
    INIT => X"0080"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA_1_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(5),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xzAregLoadEn_1: LUT2 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2023,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_1);
  x_g0_rn: LUT4 
  generic map(
    INIT => X"0E0A"
  )
  port map (
    I0 => G2_4,
    I1 => G4_5,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(57),
    O => G0_RN_0);
  x_g0_sn: LUT4 
  generic map(
    INIT => X"0040"
  )
  port map (
    I0 => G2_4,
    I1 => G4_5,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    O => G0_SN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_sqmuxa_1_1: LUT4 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => N_12791,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(5),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_25_0_0: LUT4 
  generic map(
    INIT => X"E33C"
  )
  port map (
    I0 => N_12941,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_25_0_0_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(48),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(51),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_371);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_9_sqmuxa_m1_e_1: LUT3 
  generic map(
    INIT => X"7F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA_M1_E_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(5),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA_M1_E_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_9_sqmuxa_m1_e: LUT4 
  generic map(
    INIT => X"0E02"
  )
  port map (
    I0 => G0_RN_0,
    I1 => G0_SN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA_M1_E_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(57),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_3_1: LUT2 
  generic map(
    INIT => X"6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_3_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_expaddershft_un42_expxbus_3: LUT4_L 
  generic map(
    INIT => X"E12D"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_853,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_854,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_3_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_m5_0x: LUT3 
  generic map(
    INIT => X"F2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M14(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_0X(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_2_0_rn_3x: LUT3 
  generic map(
    INIT => X"5C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2017,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(241),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_0_RN_0(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_2_0_3x: LUT3 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_0_RN_0(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_0X(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_853);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m14_0_amx_3x: LUT4 
  generic map(
    INIT => X"0002"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_53_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(8),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(9),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M14_0X(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m14_0_bmx_3x: LUT4 
  generic map(
    INIT => X"F7FF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SM0_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SM3_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV_4_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M14_0X_0(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_21_i_L5: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(41),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(42),
    O => N_12973);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_23_i_L5: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(43),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(44),
    O => N_13005);
  x_g0_L1: LUT3 
  generic map(
    INIT => X"15"
  )
  port map (
    I0 => G2_4,
    I1 => G4_5,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(57),
    O => N_13009);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_28_0_sn: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(49),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(50),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_18_0_0x: LUT4_L 
  generic map(
    INIT => X"ACA3"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_363,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(51),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(52),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_26_0_0X);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_26_0_0_rn_1: LUT2 
  generic map(
    INIT => X"6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_25_0_0_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(48),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_26_0_0_RN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_26_0_0_rn: LUT4_L 
  generic map(
    INIT => X"5CAC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_26_0_0_RN_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_26_0_0X,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(50),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(51),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_26_0_0_RN_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_26_0_0_sn: LUT4 
  generic map(
    INIT => X"4000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_25_0_0_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(48),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(50),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(51),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_26_0_0_SN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_26_0_0: LUT3_L 
  generic map(
    INIT => X"AC"
  )
  port map (
    I0 => N_12941,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_26_0_0_RN_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_26_0_0_SN,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_372);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_1_2x: LUT2 
  generic map(
    INIT => X"7"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(10),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS_0_0_0_1(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_2x: LUT4 
  generic map(
    INIT => X"E4CC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(54),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(229),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS_0_0_0_1(5),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_109);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_2_L1: LUT2_L 
  generic map(
    INIT => X"6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    LO => N_13011);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_3x: LUT4 
  generic map(
    INIT => X"E4CC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(228),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS_0_0_0_1(5),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_110);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_6_sqmuxa_1: LUT2 
  generic map(
    INIT => X"7"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA_1_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_6_sqmuxa: LUT4 
  generic map(
    INIT => X"0002"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(5),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_47_i_L15: LUT3 
  generic map(
    INIT => X"53"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    O => N_13062);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_47_i_L13: LUT3_L 
  generic map(
    INIT => X"45"
  )
  port map (
    I0 => N_13060,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    LO => N_13061);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_47_i_L11: LUT4_L 
  generic map(
    INIT => X"ECA0"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(7),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(50),
    LO => N_13060);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_51_i_L14: LUT4 
  generic map(
    INIT => X"53FF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(10),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    O => N_13088);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_53_i_L14: LUT4 
  generic map(
    INIT => X"53FF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(12),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(14),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    O => N_13113);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_notsrres_m_1_1_57x: LUT3 
  generic map(
    INIT => X"08"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_FPLD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA_1_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(5),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_1_1(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_notsrres_m_1_57x: LUT4 
  generic map(
    INIT => X"0040"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_1_1(57),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_1(57));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_6_i_L1: LUT2_L 
  generic map(
    INIT => X"7"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_6_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_6_6,
    LO => N_13133);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_7_sqmuxa: LUT4 
  generic map(
    INIT => X"8000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_1_1(57),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_24_i_L1: LUT4 
  generic map(
    INIT => X"040C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_24_4,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M_0(44),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(45),
    O => N_13154);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_48_i_L1: LUT4 
  generic map(
    INIT => X"040C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_48_4,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M_0(8),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(9),
    O => N_13175);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_52_i_L1: LUT4 
  generic map(
    INIT => X"040C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_52_4,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M_0(12),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(13),
    O => N_13196);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_22_i_L1: LUT4 
  generic map(
    INIT => X"040C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_22_4,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M_0(42),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(43),
    O => N_13217);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_54_i_L1: LUT4 
  generic map(
    INIT => X"040C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_54_4,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M_0(14),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(15),
    O => N_13238);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_8_sqmuxa: LUT4 
  generic map(
    INIT => X"4000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_1_1(57),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_m_0_1_3x: LUT4 
  generic map(
    INIT => X"5506"
  )
  port map (
    I0 => N_12614,
    I1 => N_12615,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_M_0_1(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_4x: LUT4 
  generic map(
    INIT => X"E4CC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(52),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(227),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS_0_0_0_1(5),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_111);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_c_fax_xzybus_0_0_0_5x: LUT4 
  generic map(
    INIT => X"E4CC"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(226),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS_0_0_0_1(5),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_112);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_28_0_rn_0: LUT4 
  generic map(
    INIT => X"1CC3"
  )
  port map (
    I0 => N_12941,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_25_0_0_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(48),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(51),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_28_0: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1519);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_m_0_1_5x: LUT4 
  generic map(
    INIT => X"0E1F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT0(5),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(5),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_M_0_1(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_m_0_1_6x: LUT4 
  generic map(
    INIT => X"0E1F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT0(6),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(6),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_M_0_1(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_m_0_1_7x: LUT4 
  generic map(
    INIT => X"0E1F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT0(7),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_M_0_1(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_m_0_1_1x: LUT4 
  generic map(
    INIT => X"0E1F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT0(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_M_0_1(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_m_0_1_0x: LUT4 
  generic map(
    INIT => X"0E1F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT0(0),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_M_0_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_m_0_1_2x: LUT4 
  generic map(
    INIT => X"0E1F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT0(2),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_M_0_1(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_m_0_L1: LUT4 
  generic map(
    INIT => X"0E1F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT0(4),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(4),
    O => N_13323);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_25_0_0_L9_L3: LUT3 
  generic map(
    INIT => X"7F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(51),
    I1 => GRLFPC2_0_FPO_FRAC(52),
    I2 => GRLFPC2_0_FPO_FRAC(53),
    O => N_13349);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_wqstsets_1_0_9x: LUT4 
  generic map(
    INIT => X"028A"
  )
  port map (
    I0 => N_13359,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(56),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_WQSTSETS_1_0(9));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_wqstsets_1_0_L1: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(55),
    O => N_13359);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xzBregLoadEn_1: LUT4_L 
  generic map(
    INIT => X"111A"
  )
  port map (
    I0 => G0_SN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(3),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xzBregLoadEn: LUT4 
  generic map(
    INIT => X"1C10"
  )
  port map (
    I0 => N_13009,
    I1 => G0_SN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(57),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZBREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_2_m_0_1_8x: LUT4 
  generic map(
    INIT => X"5F3F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M_0_1(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_2_m_0_8x: LUT4 
  generic map(
    INIT => X"0080"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_1_1(57),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M_0_1(8),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M_0(8));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_2_m_0_1_14x: LUT4 
  generic map(
    INIT => X"5F3F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(12),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(14),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M_0_1(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_2_m_0_14x: LUT4 
  generic map(
    INIT => X"0080"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_1_1(57),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M_0_1(14),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M_0(14));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_2_m_0_1_42x: LUT4 
  generic map(
    INIT => X"5F3F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(40),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M_0_1(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_2_m_0_42x: LUT4 
  generic map(
    INIT => X"0080"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_1_1(57),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M_0_1(42),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M_0(42));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_2_m_0_1_12x: LUT4 
  generic map(
    INIT => X"5F3F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(10),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M_0_1(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_2_m_0_12x: LUT4 
  generic map(
    INIT => X"0080"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_1_1(57),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M_0_1(12),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M_0(12));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_2_m_0_1_44x: LUT4 
  generic map(
    INIT => X"5F3F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(42),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_4(44),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M_0_1(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_s_1_2_m_0_44x: LUT4 
  generic map(
    INIT => X"0080"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_1_1(57),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M_0_1(44),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M_0(44));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_countsuccessivezero_m12_0_0x: LUT4_L 
  generic map(
    INIT => X"CAAA"
  )
  port map (
    I0 => N_12106,
    I1 => N_12107,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_53_I,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV_6_1,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M12(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_r_dpath_inv_6_1_0: LUT2 
  generic map(
    INIT => X"1"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(4),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(6),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV_6_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_r_dpath_inv_6: LUT4 
  generic map(
    INIT => X"1000"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV_6_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV_6_1_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_25_0_0_L9_L7_1: LUT3 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(56),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(56),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_25_0_0_L9_L7_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_sqmuxa_1_1_0: LUT3_L 
  generic map(
    INIT => X"1B"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(57),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(57),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_1_sqmuxa_1: LUT4 
  generic map(
    INIT => X"0A0E"
  )
  port map (
    I0 => G2_4,
    I1 => G4_5,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1_1_0,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_SQMUXA_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_53_i_1: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(13),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(14),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_53_I_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_51_i_1: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(11),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(12),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_51_I_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_1_176x: LUT3 
  generic map(
    INIT => X"68"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTXZYFROMD_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_0_1(176));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_0_0_176x: LUT3 
  generic map(
    INIT => X"E4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_0_1(176),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(55),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_278);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_2_1_1_0_1x: LUT4_L 
  generic map(
    INIT => X"2FAF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_I_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(10),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_2_1_1_0(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_xzybus_2_1_1x: LUT4_L 
  generic map(
    INIT => X"4044"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN5_XZYBUSLSBS,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_2_1_1_0(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTXZYFROMD_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(230),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_2_1(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_fast_375x: FDS port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_FAST(375),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_1_I(375),
      C => clk,
      S => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_0_I(375));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un4_notxzyfromd_i_sx: LUT4_L 
  generic map(
    INIT => X"EAC0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_DREG_FAST(51),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_FAST(376),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(9),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(14),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_I_SX);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un4_notxzyfromd_i: LUT3 
  generic map(
    INIT => X"15"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN4_NOTXZYFROMD_I_SX,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(10),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2263_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_6_1: LUT2 
  generic map(
    INIT => X"6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_6_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_feedback_0_0x: LUT4 
  generic map(
    INIT => X"1F10"
  )
  port map (
    I0 => N_2477,
    I1 => N_13799,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACKMULXFF_UN18_FEEDBACK,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(60),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_FEEDBACK(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_feedback_0_L1: LUT4_L 
  generic map(
    INIT => X"1051"
  )
  port map (
    I0 => N_2476,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN20_LOCOV_5,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN30_LOCOV_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    LO => N_13799);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_rn_2x: LUT4 
  generic map(
    INIT => X"2320"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_846,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_854,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_RN_0(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_sn_2x: LUT4 
  generic map(
    INIT => X"0001"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_854,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_SN(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_2x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_RN_0(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_SN(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M14(2),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_rn_1x: LUT4 
  generic map(
    INIT => X"2320"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_845,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_854,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_RN_1(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_sn_1x: LUT4 
  generic map(
    INIT => X"0001"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_854,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_SN(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_1x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_RN_1(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_SN(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M14(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_0_L3: LUT4_L 
  generic map(
    INIT => X"0C0A"
  )
  port map (
    I0 => N_12164,
    I1 => N_12165,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(2),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV_6,
    LO => N_14071);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_rn_0x: LUT4 
  generic map(
    INIT => X"2320"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_844,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_854,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_RN_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_sn_0x: LUT4 
  generic map(
    INIT => X"0001"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_854,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_SN(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_0x: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_RN_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_SN(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_M14(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_dpath_new_8_sqmuxa_1_1: LUT3 
  generic map(
    INIT => X"40"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2023,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(7),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA_1_1);
  x_g0_L1_0: LUT3 
  generic map(
    INIT => X"15"
  )
  port map (
    I0 => G2_4,
    I1 => G4_5,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(57),
    O => N_14297);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_r_dpath_inv: LUT4 
  generic map(
    INIT => X"4000"
  )
  port map (
    I0 => N_14349,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_53_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_COUNTSUCCESSIVEZERO_SM3_I,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV_6_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_r_dpath_inv_L1: LUT4_L 
  generic map(
    INIT => X"0001"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(15),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(16),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(17),
    LO => N_14348);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_25_0_0_L9_L1_1: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(47),
    I1 => GRLFPC2_0_FPO_FRAC(48),
    I2 => GRLFPC2_0_FPO_FRAC(49),
    I3 => GRLFPC2_0_FPO_FRAC(50),
    LO => N_14411);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_28_0_rn_rn_1: LUT2 
  generic map(
    INIT => X"6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZZERO_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(52),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_RN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_28_0_rn_1: LUT3_L 
  generic map(
    INIT => X"5C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_363,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_RN_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(51),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_28_0_rn: LUT4 
  generic map(
    INIT => X"C044"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_361,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_1_0,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(49),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_0_1_0_3x: LUT4_L 
  generic map(
    INIT => X"3035"
  )
  port map (
    I0 => N_14071,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_847,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_R_DPATH_INV,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_1_0(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_leftshifterbl_slcontrol_0_3x: LUT3 
  generic map(
    INIT => X"B1"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_854,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_1_0(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m3_0_sx: LUT4_L 
  generic map(
    INIT => X"4FEF"
  )
  port map (
    I0 => G0_SN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(3),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(57),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_M3_0_SX);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_rin_dpath_sn_m3_0: LUT3 
  generic map(
    INIT => X"0D"
  )
  port map (
    I0 => N_14297,
    I1 => G0_SN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH_SN_M3_0_SX,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_740);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un21_notxzyfromd_i_sx: LUT4_L 
  generic map(
    INIT => X"F888"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_DREG_FAST(53),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_FAST(375),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(11),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(13),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_I_SX);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_fax_un21_notxzyfromd_i: LUT3 
  generic map(
    INIT => X"45"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN21_NOTXZYFROMD_I_SX,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(10),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_25_0_0_L9_L1_L1: LUT3 
  generic map(
    INIT => X"01"
  )
  port map (
    I0 => N_2476,
    I1 => N_2477,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_UN42_EXPXBUS,
    O => N_15046);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_25_0_0_L9: LUT4 
  generic map(
    INIT => X"8CC0"
  )
  port map (
    I0 => N_13349,
    I1 => N_15069,
    I2 => N_15070,
    I3 => GRLFPC2_0_FPO_FRAC(54),
    O => N_12941);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_25_0_0_L9_L3_1: LUT4_L 
  generic map(
    INIT => X"353F"
  )
  port map (
    I0 => N_13359,
    I1 => N_14411,
    I2 => GRLFPC2_0_FPO_FRAC(54),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_25_0_0_L9_L7_1,
    LO => N_15070);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_notsqrtlftcc_1_25_0_0_L9_L1_2: LUT4 
  generic map(
    INIT => X"20A2"
  )
  port map (
    I0 => N_15046,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN20_LOCOV_5,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_REEXCOVUV_UN30_LOCOV_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0,
    O => N_15069);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un4_temp_2_0_rn_0x: LUT3 
  generic map(
    INIT => X"D8"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(24),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(25),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN4_TEMP_2_0_RN_1(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un4_temp_2_0_0x: LUT3 
  generic map(
    INIT => X"CA"
  )
  port map (
    I0 => N_12084,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN4_TEMP_2_0_RN_1(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_UN1_GRFPULITE0_FAST,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_104);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xzAregLoadEn_rn: LUT4_L 
  generic map(
    INIT => X"E0A0"
  )
  port map (
    I0 => G2_4,
    I1 => G4_5,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(57),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_RN_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xzAregLoadEn_sn: LUT4 
  generic map(
    INIT => X"4000"
  )
  port map (
    I0 => G2_4,
    I1 => G4_5,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_SN_N_4,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_SN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_dpxx_xzAregLoadEn: LUT3 
  generic map(
    INIT => X"E2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_RN_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN_SN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(57),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_21_i_1_0: LUT4_L 
  generic map(
    INIT => X"40C0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_21_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_21_4,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(42),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_21_I_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_23_i_1_0: LUT4_L 
  generic map(
    INIT => X"40C0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_23_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_23_4,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(44),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_23_I_1_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_47_i_L3: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => N_13062,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_0(8),
    O => N_15368);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_47_i_L1_0: LUT3 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN1_XZYBUS24_S0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_47_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(8),
    O => N_15367);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_51_i_L10: LUT4_L 
  generic map(
    INIT => X"FDDD"
  )
  port map (
    I0 => N_15387,
    I1 => N_15388,
    I2 => N_15389,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    LO => N_13086);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_51_i_L10_L15: LUT4 
  generic map(
    INIT => X"5044"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(13),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => N_15389);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_51_i_L10_L13: LUT3_L 
  generic map(
    INIT => X"D5"
  )
  port map (
    I0 => N_15386,
    I1 => GRLFPC2_0_FPO_FRAC(11),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    LO => N_15388);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_51_i_L10_L10: LUT2 
  generic map(
    INIT => X"7"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(46),
    O => N_15387);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_51_i_L10_L6: LUT3 
  generic map(
    INIT => X"15"
  )
  port map (
    I0 => N_15385,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(45),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    O => N_15386);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_51_i_L10_L4: LUT4_L 
  generic map(
    INIT => X"DC50"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(45),
    I3 => rfo2_data2(9),
    LO => N_15385);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_53_i_L10: LUT4_L 
  generic map(
    INIT => X"FDDD"
  )
  port map (
    I0 => N_15408,
    I1 => N_15409,
    I2 => N_15410,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    LO => N_13111);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_53_i_L10_L15: LUT4 
  generic map(
    INIT => X"5044"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(14),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(15),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_WQSCTRL,
    O => N_15410);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_53_i_L10_L13: LUT3_L 
  generic map(
    INIT => X"D5"
  )
  port map (
    I0 => N_15407,
    I1 => GRLFPC2_0_FPO_FRAC(13),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    LO => N_15409);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_53_i_L10_L10: LUT2 
  generic map(
    INIT => X"7"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_3_SQMUXA_2,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(44),
    O => N_15408);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_53_i_L10_L6: LUT3 
  generic map(
    INIT => X"15"
  )
  port map (
    I0 => N_15406,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(43),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_9_SQMUXA,
    O => N_15407);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_53_i_L10_L4: LUT4_L 
  generic map(
    INIT => X"DC50"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_1_M_1(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(43),
    I3 => rfo2_data2(11),
    LO => N_15406);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_30_i_L8: LUT4_L 
  generic map(
    INIT => X"1300"
  )
  port map (
    I0 => N_15500,
    I1 => N_15501,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_30_0,
    LO => N_15502);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_30_i_L6: LUT2 
  generic map(
    INIT => X"4"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZAREGLOADEN,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(36),
    O => N_15501);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_30_i_L4: LUT3 
  generic map(
    INIT => X"01"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRTOSTICKY_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_SE(21),
    O => N_15500);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_6_i_1: LUT4 
  generic map(
    INIT => X"4C5F"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(52),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(52),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_6_I_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_5_i_L3: LUT4_L 
  generic map(
    INIT => X"048C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SRCONTROL_1(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_1(57),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(52),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_2(53),
    LO => N_15543);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_55_i_1: LUT4 
  generic map(
    INIT => X"00B0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_6_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_55_0,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0_M(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_55_I_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_8_i_L5: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(55),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(59),
    O => N_15777);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_8_i_L3: LUT2 
  generic map(
    INIT => X"7"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_278,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    O => N_15776);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_8_i_L1: LUT4 
  generic map(
    INIT => X"40C0"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_1(57),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_8_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_8_5,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(56),
    O => N_15775);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_7_i_L8: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(53),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(61),
    O => N_15809);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_7_i_L6: LUT4_L 
  generic map(
    INIT => X"BF3F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_1(57),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_7_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_7_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(54),
    LO => N_15808);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_7_i_L3: LUT2 
  generic map(
    INIT => X"7"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(53),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    O => N_15807);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_2_i_L8: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(48),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
    O => N_15822);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_2_i_L6: LUT4_L 
  generic map(
    INIT => X"BF3F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_1(57),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_2_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_2_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(49),
    LO => N_15821);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_2_i_L3: LUT2 
  generic map(
    INIT => X"7"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(48),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    O => N_15820);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_1_i_L8: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(47),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(67),
    O => N_15854);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_1_i_L6: LUT4_L 
  generic map(
    INIT => X"BF3F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_1(57),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_1_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_1_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(48),
    LO => N_15853);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_1_i_L3: LUT2 
  generic map(
    INIT => X"7"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(47),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    O => N_15852);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_3_i_L5: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(49),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(65),
    O => N_15885);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_3_i_L3: LUT4 
  generic map(
    INIT => X"0700"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(49),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH_M(7),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_3_0,
    O => N_15884);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_3_i_L1: LUT3 
  generic map(
    INIT => X"4C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_1(57),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_3_6,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(50),
    O => N_15883);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_4_i_L8: LUT4 
  generic map(
    INIT => X"23AF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(50),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_2_SQMUXA_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
    O => N_15898);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_4_i_L6: LUT4_L 
  generic map(
    INIT => X"BF3F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_1(57),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_4_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_4_6,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1(51),
    LO => N_15897);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_4_i_L3: LUT2 
  generic map(
    INIT => X"7"
  )
  port map (
    I0 => GRLFPC2_0_FPO_FRAC(50),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    O => N_15896);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_9_i_1: LUT4 
  generic map(
    INIT => X"4FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_RIGHTSHIFTERBL_S_8(57),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M_1(57),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_9_0,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_9_5,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_9_I_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_5_i_1: LUT4_L 
  generic map(
    INIT => X"1500"
  )
  port map (
    I0 => N_15543,
    I1 => GRLFPC2_0_FPO_FRAC(51),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_5_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_5_6,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_5_I_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_30_i_1: LUT3_L 
  generic map(
    INIT => X"75"
  )
  port map (
    I0 => N_15502,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(20),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_7_SQMUXA,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_30_I_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_7_1: LUT2 
  generic map(
    INIT => X"6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(7),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_7_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_8_1: LUT2 
  generic map(
    INIT => X"6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(8),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_8_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_9_1: LUT2 
  generic map(
    INIT => X"6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(9),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_9_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_10_1: LUT2 
  generic map(
    INIT => X"6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(10),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_10_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_11_1: LUT2 
  generic map(
    INIT => X"6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(11),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_11_1);
  x_g0: LUT4 
  generic map(
    INIT => X"CD01"
  )
  port map (
    I0 => N_20103,
    I1 => G0_SN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF1(57),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_SXC_SFTLFT_UN4_AREGSIGN_SEL);
  x_g0_L1_1: LUT3_L 
  generic map(
    INIT => X"15"
  )
  port map (
    I0 => G2_4,
    I1 => G4_5,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUF0(57),
    LO => N_20103);
  x_grlfpc2_0_r_mk_rstc_1_0: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => GRLFPC2_0_N_782,
    I1 => GRLFPC2_0_R_MK_HOLDN2,
    I2 => GRLFPC2_0_R_MK_HOLDN1,
    O => GRLFPC2_0_R_MK_RSTC_1_0);
  x_grlfpc2_0_comb_fpdecode_un1_wren210_2: LUT3 
  generic map(
    INIT => X"08"
  )
  port map (
    I0 => GRLFPC2_0_MOV_2_SQMUXA_1_0,
    I1 => cpi_d_inst(11),
    I2 => cpi_d_inst(10),
    O => GRLFPC2_0_COMB_FPDECODE_RS2D5_3);
  x_grlfpc2_0_rs2_0_sqmuxa: LUT3 
  generic map(
    INIT => X"08"
  )
  port map (
    I0 => GRLFPC2_0_COMB_FPDECODE_UN3_OP,
    I1 => cpi_d_inst(31),
    I2 => cpi_d_inst(30),
    O => GRLFPC2_0_RS2_0_SQMUXA);
  x_grlfpc2_0_rs1v_1_sqmuxa: LUT3 
  generic map(
    INIT => X"04"
  )
  port map (
    I0 => GRLFPC2_0_COMB_FPDECODE_MOV11,
    I1 => cpi_d_inst(31),
    I2 => cpi_d_inst(30),
    O => GRLFPC2_0_RS1V_1_SQMUXA);
  x_grlfpc2_0_rs1v_0_sqmuxa: LUT3 
  generic map(
    INIT => X"40"
  )
  port map (
    I0 => GRLFPC2_0_RS1V10_I,
    I1 => cpi_d_inst(31),
    I2 => cpi_d_inst(30),
    O => GRLFPC2_0_RS1V_0_SQMUXA);
  x_grlfpc2_0_comb_v_e_stdata_1_1_bm_0x: LUT3 
  generic map(
    INIT => X"8A"
  )
  port map (
    I0 => GRLFPC2_0_R_I_INST(0),
    I1 => cpi_a_cnt(1),
    I2 => cpi_a_cnt(0),
    O => N_12219);
  x_grlfpc2_0_comb_v_e_stdata_1_2_bm_1x: LUT3 
  generic map(
    INIT => X"8A"
  )
  port map (
    I0 => GRLFPC2_0_R_I_INST(1),
    I1 => cpi_a_cnt(1),
    I2 => cpi_a_cnt(0),
    O => N_12257);
  x_grlfpc2_0_wren1_1_sqmuxa_1: LUT3 
  generic map(
    INIT => X"02"
  )
  port map (
    I0 => GRLFPC2_0_WREN2_1_SQMUXA_1_0,
    I1 => cpi_x_cnt(1),
    I2 => cpi_x_cnt(0),
    O => GRLFPC2_0_WREN1_1_SQMUXA_1);
  x_grlfpc2_0_wraddr_0_sqmuxa: LUT3 
  generic map(
    INIT => X"40"
  )
  port map (
    I0 => cpi_dbg_fsr,
    I1 => cpi_dbg_write,
    I2 => cpi_dbg_enable,
    O => GRLFPC2_0_WRADDR_0_SQMUXA);
  x_grlfpc2_0_v_fsr_nonstd_0_sqmuxa_1: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => cpi_dbg_fsr,
    I1 => cpi_dbg_write,
    I2 => cpi_dbg_enable,
    O => GRLFPC2_0_V_FSR_NONSTD_0_SQMUXA_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_r_dpath_inv_L3: LUT3_L 
  generic map(
    INIT => X"FD"
  )
  port map (
    I0 => N_14348,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(14),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(13),
    LO => N_14349);
  x_grlfpc2_0_un1_holdn_1: LUT3 
  generic map(
    INIT => X"15"
  )
  port map (
    I0 => GRLFPC2_0_COMB_UN6_IUEXEC,
    I1 => holdn,
    I2 => GRLFPC2_0_N_691,
    O => GRLFPC2_0_N_762);
  x_grlfpc2_0_I_205: LUT3 
  generic map(
    INIT => X"80"
  )
  port map (
    I0 => cpi_d_inst(0),
    I1 => GRLFPC2_0_MOV_7_SQMUXA_3,
    I2 => cpi_d_inst(23),
    O => GRLFPC2_0_N_654);
  x_grlfpc2_0_comb_fpdecode_mov11: LUT3 
  generic map(
    INIT => X"40"
  )
  port map (
    I0 => cpi_d_inst(19),
    I1 => GRLFPC2_0_MOV_7_SQMUXA_3,
    I2 => cpi_d_inst(23),
    O => GRLFPC2_0_COMB_FPDECODE_MOV11);
  x_grlfpc2_0_un1_afq3: LUT3 
  generic map(
    INIT => X"5D"
  )
  port map (
    I0 => GRLFPC2_0_COMB_FPDECODE_AFQ4_1,
    I1 => cpi_d_inst(20),
    I2 => cpi_d_inst(19),
    O => GRLFPC2_0_UN1_AFQ3_I);
  x_grlfpc2_0_N_762_i: LUT3 
  generic map(
    INIT => X"F8"
  )
  port map (
    I0 => GRLFPC2_0_N_691,
    I1 => holdn,
    I2 => GRLFPC2_0_COMB_UN6_IUEXEC,
    O => GRLFPC2_0_N_762_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_fast_53x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_DREG_FAST(53),
      D => N_6882_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_45_rep2: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
      D => N_6874_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_45_rep1: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
      D => N_6874_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_fast_45x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_FAST(17),
      D => N_6874_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_46_rep1: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_16_REP1,
      D => N_6875_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_fast_46x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_FAST(16),
      D => N_6875_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_fast_51x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_DREG_FAST(51),
      D => N_6880_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_r_x_seqerr_0_0_DOUT_0x: FDE port map (
      Q => GRLFPC2_0_R_X_SEQERR,
      D => GRLFPC2_0_R_X_SEQERR_0_0_N_6,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_x_rdd_0_0_DOUT_0x: FDE port map (
      Q => GRLFPC2_0_R_X_RDD,
      D => GRLFPC2_0_R_X_RDD_0_0_TMP_D_ARRAY_0(0),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_areg_1x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(1),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_REP1,
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_areg_0x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(0),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_0_REP1,
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_areg_7x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(7),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_6_REP1,
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_areg_6x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(6),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_5_REP1,
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_areg_5x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(5),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_3_REP1,
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_areg_4x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(4),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_2_REP1,
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_areg_3x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(3),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_7_REP1,
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_areg_2x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_PCTRL_NEW_19_0_AREG(2),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_4_REP1,
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_62x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(0),
      D => N_6891_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_61x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(1),
      D => N_6890_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_60x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(2),
      D => N_6889_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_59x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(3),
      D => N_6888_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_58x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(4),
      D => N_6887_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_57x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(5),
      D => N_6886_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_56x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(6),
      D => N_6885_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_55x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(7),
      D => N_6884_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_54x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(8),
      D => N_6883_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_53x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(9),
      D => N_6882_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_52x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(10),
      D => N_6881_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_51x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(11),
      D => N_6880_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_50x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(12),
      D => N_6879_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_49x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(13),
      D => N_6878_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_48x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(14),
      D => N_6877_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_47x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_I(15),
      D => N_6876_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_46x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(16),
      D => N_6875_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_45x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
      D => N_6874_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_44x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(18),
      D => N_6873_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_43x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_I(19),
      D => N_6872_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_42x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(20),
      D => N_6871_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_41x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(21),
      D => N_6870_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_40x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_I(22),
      D => N_6869_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_39x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(23),
      D => N_6868_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_38x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_I(24),
      D => N_6867_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_37x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(25),
      D => N_6866_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_36x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(26),
      D => N_6865_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_35x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(27),
      D => N_6864_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_34x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(28),
      D => N_6863_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_33x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(29),
      D => N_6862_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_32x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(30),
      D => N_6861_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_31x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
      D => N_6860_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_30x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(32),
      D => N_6859_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_29x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33),
      D => N_6858_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_28x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(34),
      D => N_6857_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_27x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(35),
      D => N_6856_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_26x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
      D => N_6855_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_25x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(38),
      D => N_6854_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_24x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(39),
      D => N_6853_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_23x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(40),
      D => N_6852_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_22x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_I(41),
      D => N_6851_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_21x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(42),
      D => N_6850_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_20x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_I(43),
      D => N_6849_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_19x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(44),
      D => N_6848_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_18x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(45),
      D => N_6847_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_17x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(46),
      D => N_6846_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_16x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(47),
      D => N_6845_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_15x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(48),
      D => N_6844_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_14x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(49),
      D => N_6843_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_13x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(50),
      D => N_6842_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_12x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(51),
      D => N_6841_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_11x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(52),
      D => N_6840_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_10x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(53),
      D => N_6839_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_9x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(54),
      D => N_6838_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_8x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(55),
      D => N_6837_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_7x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(56),
      D => N_6836_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_6x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(57),
      D => N_6835_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_5x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(58),
      D => N_6834_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_4x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(59),
      D => N_6833_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_3x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(60),
      D => N_6832_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_2x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(61),
      D => N_6831_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_1x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(62),
      D => N_6830_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_pctrl_new_19_0_dreg_0x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(63),
      D => N_6829_A,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UPDATE_1);
  x_grlfpc2_0_r_mk_holdn2: FD port map (
      Q => GRLFPC2_0_R_MK_HOLDN2,
      D => GRLFPC2_0_R_MK_HOLDN1,
      C => clk);
  x_grlfpc2_0_r_mk_rst2: FD port map (
      Q => GRLFPC2_0_R_MK_RST2,
      D => GRLFPC2_0_R_MK_RST,
      C => clk);
  x_grlfpc2_0_r_i_res_1x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(1),
      D => GRLFPC2_0_FPO_FRAC(4),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_0x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(0),
      D => GRLFPC2_0_FPO_FRAC(3),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_a_rs1_4x: FD port map (
      Q => GRLFPC2_0_R_A_RS1(4),
      D => GRLFPC2_0_COMB_RS1_1(4),
      C => clk);
  x_grlfpc2_0_r_a_rs1_3x: FD port map (
      Q => GRLFPC2_0_R_A_RS1(3),
      D => GRLFPC2_0_COMB_RS1_1(3),
      C => clk);
  x_grlfpc2_0_r_a_rs1_2x: FD port map (
      Q => GRLFPC2_0_R_A_RS1(2),
      D => GRLFPC2_0_COMB_RS1_1(2),
      C => clk);
  x_grlfpc2_0_r_a_rs1_1x: FD port map (
      Q => GRLFPC2_0_R_A_RS1(1),
      D => GRLFPC2_0_COMB_RS1_1(1),
      C => clk);
  x_grlfpc2_0_r_a_rs1_0x: FD port map (
      Q => GRLFPC2_0_R_A_RS1(0),
      D => GRLFPC2_0_COMB_RS1_1(0),
      C => clk);
  x_grlfpc2_0_r_i_res_16x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(16),
      D => GRLFPC2_0_FPO_FRAC(19),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_15x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(15),
      D => GRLFPC2_0_FPO_FRAC(18),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_14x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(14),
      D => GRLFPC2_0_FPO_FRAC(17),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_13x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(13),
      D => GRLFPC2_0_FPO_FRAC(16),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_12x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(12),
      D => GRLFPC2_0_FPO_FRAC(15),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_11x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(11),
      D => GRLFPC2_0_FPO_FRAC(14),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_10x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(10),
      D => GRLFPC2_0_FPO_FRAC(13),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_9x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(9),
      D => GRLFPC2_0_FPO_FRAC(12),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_8x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(8),
      D => GRLFPC2_0_FPO_FRAC(11),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_7x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(7),
      D => GRLFPC2_0_FPO_FRAC(10),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_6x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(6),
      D => GRLFPC2_0_FPO_FRAC(9),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_5x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(5),
      D => GRLFPC2_0_FPO_FRAC(8),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_4x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(4),
      D => GRLFPC2_0_FPO_FRAC(7),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_3x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(3),
      D => GRLFPC2_0_FPO_FRAC(6),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_2x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(2),
      D => GRLFPC2_0_FPO_FRAC(5),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_31x: FD port map (
      Q => GRLFPC2_0_R_I_RES(31),
      D => GRLFPC2_0_COMB_V_I_RES_1(31),
      C => clk);
  x_grlfpc2_0_r_i_res_30x: FD port map (
      Q => GRLFPC2_0_R_I_RES(30),
      D => GRLFPC2_0_COMB_V_I_RES_1(30),
      C => clk);
  x_grlfpc2_0_r_i_res_29x: FD port map (
      Q => GRLFPC2_0_R_I_RES(29),
      D => GRLFPC2_0_COMB_V_I_RES_1(29),
      C => clk);
  x_grlfpc2_0_r_i_res_28x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(28),
      D => GRLFPC2_0_FPO_FRAC(31),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_27x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(27),
      D => GRLFPC2_0_FPO_FRAC(30),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_26x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(26),
      D => GRLFPC2_0_FPO_FRAC(29),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_25x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(25),
      D => GRLFPC2_0_FPO_FRAC(28),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_24x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(24),
      D => GRLFPC2_0_FPO_FRAC(27),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_23x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(23),
      D => GRLFPC2_0_FPO_FRAC(26),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_22x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(22),
      D => GRLFPC2_0_FPO_FRAC(25),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_21x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(21),
      D => GRLFPC2_0_FPO_FRAC(24),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_20x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(20),
      D => GRLFPC2_0_FPO_FRAC(23),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_19x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(19),
      D => GRLFPC2_0_FPO_FRAC(22),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_18x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(18),
      D => GRLFPC2_0_FPO_FRAC(21),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_17x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(17),
      D => GRLFPC2_0_FPO_FRAC(20),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_46x: FD port map (
      Q => GRLFPC2_0_R_I_RES(46),
      D => GRLFPC2_0_COMB_V_I_RES_1(46),
      C => clk);
  x_grlfpc2_0_r_i_res_45x: FD port map (
      Q => GRLFPC2_0_R_I_RES(45),
      D => GRLFPC2_0_COMB_V_I_RES_1(45),
      C => clk);
  x_grlfpc2_0_r_i_res_44x: FD port map (
      Q => GRLFPC2_0_R_I_RES(44),
      D => GRLFPC2_0_COMB_V_I_RES_1(44),
      C => clk);
  x_grlfpc2_0_r_i_res_43x: FD port map (
      Q => GRLFPC2_0_R_I_RES(43),
      D => GRLFPC2_0_COMB_V_I_RES_1(43),
      C => clk);
  x_grlfpc2_0_r_i_res_42x: FD port map (
      Q => GRLFPC2_0_R_I_RES(42),
      D => GRLFPC2_0_COMB_V_I_RES_1(42),
      C => clk);
  x_grlfpc2_0_r_i_res_41x: FD port map (
      Q => GRLFPC2_0_R_I_RES(41),
      D => GRLFPC2_0_COMB_V_I_RES_1(41),
      C => clk);
  x_grlfpc2_0_r_i_res_40x: FD port map (
      Q => GRLFPC2_0_R_I_RES(40),
      D => GRLFPC2_0_COMB_V_I_RES_1(40),
      C => clk);
  x_grlfpc2_0_r_i_res_39x: FD port map (
      Q => GRLFPC2_0_R_I_RES(39),
      D => GRLFPC2_0_COMB_V_I_RES_1(39),
      C => clk);
  x_grlfpc2_0_r_i_res_38x: FD port map (
      Q => GRLFPC2_0_R_I_RES(38),
      D => GRLFPC2_0_COMB_V_I_RES_1(38),
      C => clk);
  x_grlfpc2_0_r_i_res_37x: FD port map (
      Q => GRLFPC2_0_R_I_RES(37),
      D => GRLFPC2_0_COMB_V_I_RES_1(37),
      C => clk);
  x_grlfpc2_0_r_i_res_36x: FD port map (
      Q => GRLFPC2_0_R_I_RES(36),
      D => GRLFPC2_0_COMB_V_I_RES_1(36),
      C => clk);
  x_grlfpc2_0_r_i_res_35x: FD port map (
      Q => GRLFPC2_0_R_I_RES(35),
      D => GRLFPC2_0_COMB_V_I_RES_1(35),
      C => clk);
  x_grlfpc2_0_r_i_res_34x: FD port map (
      Q => GRLFPC2_0_R_I_RES(34),
      D => GRLFPC2_0_COMB_V_I_RES_1(34),
      C => clk);
  x_grlfpc2_0_r_i_res_33x: FD port map (
      Q => GRLFPC2_0_R_I_RES(33),
      D => GRLFPC2_0_COMB_V_I_RES_1(33),
      C => clk);
  x_grlfpc2_0_r_i_res_32x: FD port map (
      Q => GRLFPC2_0_R_I_RES(32),
      D => GRLFPC2_0_COMB_V_I_RES_1(32),
      C => clk);
  x_grlfpc2_0_r_i_res_61x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(61),
      D => GRLFPC2_0_FPO_EXP(9),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_60x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(60),
      D => GRLFPC2_0_FPO_EXP(8),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_res_59x: FD port map (
      Q => GRLFPC2_0_R_I_RES(59),
      D => GRLFPC2_0_COMB_V_I_RES_1(59),
      C => clk);
  x_grlfpc2_0_r_i_res_58x: FD port map (
      Q => GRLFPC2_0_R_I_RES(58),
      D => GRLFPC2_0_COMB_V_I_RES_1(58),
      C => clk);
  x_grlfpc2_0_r_i_res_57x: FD port map (
      Q => GRLFPC2_0_R_I_RES(57),
      D => GRLFPC2_0_COMB_V_I_RES_1(57),
      C => clk);
  x_grlfpc2_0_r_i_res_56x: FD port map (
      Q => GRLFPC2_0_R_I_RES(56),
      D => GRLFPC2_0_COMB_V_I_RES_1(56),
      C => clk);
  x_grlfpc2_0_r_i_res_55x: FD port map (
      Q => GRLFPC2_0_R_I_RES(55),
      D => GRLFPC2_0_COMB_V_I_RES_1(55),
      C => clk);
  x_grlfpc2_0_r_i_res_54x: FD port map (
      Q => GRLFPC2_0_R_I_RES(54),
      D => GRLFPC2_0_COMB_V_I_RES_1(54),
      C => clk);
  x_grlfpc2_0_r_i_res_53x: FD port map (
      Q => GRLFPC2_0_R_I_RES(53),
      D => GRLFPC2_0_COMB_V_I_RES_1(53),
      C => clk);
  x_grlfpc2_0_r_i_res_52x: FD port map (
      Q => GRLFPC2_0_R_I_RES(52),
      D => GRLFPC2_0_COMB_V_I_RES_1(52),
      C => clk);
  x_grlfpc2_0_r_i_res_51x: FD port map (
      Q => GRLFPC2_0_R_I_RES(51),
      D => GRLFPC2_0_COMB_V_I_RES_1(51),
      C => clk);
  x_grlfpc2_0_r_i_res_50x: FD port map (
      Q => GRLFPC2_0_R_I_RES(50),
      D => GRLFPC2_0_COMB_V_I_RES_1(50),
      C => clk);
  x_grlfpc2_0_r_i_res_49x: FD port map (
      Q => GRLFPC2_0_R_I_RES(49),
      D => GRLFPC2_0_COMB_V_I_RES_1(49),
      C => clk);
  x_grlfpc2_0_r_i_res_48x: FD port map (
      Q => GRLFPC2_0_R_I_RES(48),
      D => GRLFPC2_0_COMB_V_I_RES_1(48),
      C => clk);
  x_grlfpc2_0_r_i_res_47x: FD port map (
      Q => GRLFPC2_0_R_I_RES(47),
      D => GRLFPC2_0_COMB_V_I_RES_1(47),
      C => clk);
  x_grlfpc2_0_r_i_res_63x: FD port map (
      Q => GRLFPC2_0_R_I_RES(63),
      D => GRLFPC2_0_COMB_V_I_RES_1(63),
      C => clk);
  x_grlfpc2_0_r_i_res_62x: FDE port map (
      Q => GRLFPC2_0_R_I_RES(62),
      D => GRLFPC2_0_FPO_EXP(10),
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_e_afq: FDE port map (
      Q => GRLFPC2_0_R_E_AFQ,
      D => GRLFPC2_0_COMB_V_E_AFQ_1,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_afsr: FDE port map (
      Q => GRLFPC2_0_R_E_AFSR,
      D => GRLFPC2_0_COMB_V_E_AFSR_1,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_fpop: FDE port map (
      Q => GRLFPC2_0_R_E_FPOP,
      D => GRLFPC2_0_COMB_V_E_FPOP_1,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_ld: FDE port map (
      Q => GRLFPC2_0_R_E_LD,
      D => GRLFPC2_0_COMB_V_E_LD_1,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_m_afq: FDE port map (
      Q => GRLFPC2_0_R_M_AFQ,
      D => GRLFPC2_0_COMB_V_M_AFQ_1,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_m_afsr: FDE port map (
      Q => GRLFPC2_0_R_M_AFSR,
      D => GRLFPC2_0_COMB_V_M_AFSR_1,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_m_fpop: FDE port map (
      Q => GRLFPC2_0_R_M_FPOP,
      D => GRLFPC2_0_COMB_V_M_FPOP_1,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_m_ld: FDE port map (
      Q => GRLFPC2_0_R_M_LD,
      D => GRLFPC2_0_COMB_V_M_LD_1,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_x_afq: FDE port map (
      Q => GRLFPC2_0_R_X_AFQ,
      D => GRLFPC2_0_COMB_V_X_AFQ_1,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_x_afsr: FDE port map (
      Q => GRLFPC2_0_R_X_AFSR,
      D => GRLFPC2_0_COMB_V_X_AFSR_1,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_x_fpop: FDE port map (
      Q => GRLFPC2_0_R_X_FPOP,
      D => GRLFPC2_0_COMB_V_X_FPOP_1,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_x_ld: FDE port map (
      Q => GRLFPC2_0_R_X_LD,
      D => GRLFPC2_0_COMB_V_X_LD_1,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_i_cc_1x: FDE port map (
      Q => GRLFPC2_0_R_I_CC(1),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1999_I,
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_cc_0x: FDE port map (
      Q => GRLFPC2_0_R_I_CC(0),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1998_I,
      C => clk,
      CE => GRLFPC2_0_COMB_UN6_IUEXEC);
  x_grlfpc2_0_r_i_inst_31x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(31),
      D => cpi_x_inst(31),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_30x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(30),
      D => cpi_x_inst(30),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_29x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(29),
      D => cpi_x_inst(29),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_28x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(28),
      D => cpi_x_inst(28),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_27x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(27),
      D => cpi_x_inst(27),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_26x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(26),
      D => cpi_x_inst(26),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_25x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(25),
      D => cpi_x_inst(25),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_24x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(24),
      D => cpi_x_inst(24),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_23x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(23),
      D => cpi_x_inst(23),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_22x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(22),
      D => cpi_x_inst(22),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_21x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(21),
      D => cpi_x_inst(21),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_20x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(20),
      D => cpi_x_inst(20),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_19x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(19),
      D => cpi_x_inst(19),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_18x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(18),
      D => cpi_x_inst(18),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_17x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(17),
      D => cpi_x_inst(17),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_16x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(16),
      D => cpi_x_inst(16),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_15x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(15),
      D => cpi_x_inst(15),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_14x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(14),
      D => cpi_x_inst(14),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_13x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(13),
      D => cpi_x_inst(13),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_12x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(12),
      D => cpi_x_inst(12),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_11x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(11),
      D => cpi_x_inst(11),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_10x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(10),
      D => cpi_x_inst(10),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_9x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(9),
      D => cpi_x_inst(9),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_8x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(8),
      D => cpi_x_inst(8),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_7x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(7),
      D => cpi_x_inst(7),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_6x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(6),
      D => cpi_x_inst(6),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_5x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(5),
      D => cpi_x_inst(5),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_4x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(4),
      D => cpi_x_inst(4),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_3x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(3),
      D => cpi_x_inst(3),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_2x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(2),
      D => cpi_x_inst(2),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_1x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(1),
      D => cpi_x_inst(1),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_inst_0x: FDE port map (
      Q => GRLFPC2_0_R_I_INST(0),
      D => cpi_x_inst(0),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_31x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(31),
      D => cpi_x_pc(31),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_30x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(30),
      D => cpi_x_pc(30),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_29x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(29),
      D => cpi_x_pc(29),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_28x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(28),
      D => cpi_x_pc(28),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_27x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(27),
      D => cpi_x_pc(27),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_26x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(26),
      D => cpi_x_pc(26),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_25x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(25),
      D => cpi_x_pc(25),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_24x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(24),
      D => cpi_x_pc(24),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_23x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(23),
      D => cpi_x_pc(23),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_22x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(22),
      D => cpi_x_pc(22),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_21x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(21),
      D => cpi_x_pc(21),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_20x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(20),
      D => cpi_x_pc(20),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_19x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(19),
      D => cpi_x_pc(19),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_18x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(18),
      D => cpi_x_pc(18),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_17x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(17),
      D => cpi_x_pc(17),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_16x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(16),
      D => cpi_x_pc(16),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_15x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(15),
      D => cpi_x_pc(15),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_14x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(14),
      D => cpi_x_pc(14),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_13x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(13),
      D => cpi_x_pc(13),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_12x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(12),
      D => cpi_x_pc(12),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_11x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(11),
      D => cpi_x_pc(11),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_10x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(10),
      D => cpi_x_pc(10),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_9x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(9),
      D => cpi_x_pc(9),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_8x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(8),
      D => cpi_x_pc(8),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_7x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(7),
      D => cpi_x_pc(7),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_6x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(6),
      D => cpi_x_pc(6),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_5x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(5),
      D => cpi_x_pc(5),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_4x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(4),
      D => cpi_x_pc(4),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_3x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(3),
      D => cpi_x_pc(3),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_i_pc_2x: FDE port map (
      Q => GRLFPC2_0_R_I_PC(2),
      D => cpi_x_pc(2),
      C => clk,
      CE => N_5258);
  x_grlfpc2_0_r_a_mov: FDE port map (
      Q => GRLFPC2_0_R_A_MOV,
      D => GRLFPC2_0_MOV_5_SQMUXA,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_i_rdd: FDE port map (
      Q => GRLFPC2_0_R_I_RDD,
      D => GRLFPC2_0_N_692,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_31x: FDE port map (
      Q => cpo_data(31),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(31),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_30x: FDE port map (
      Q => cpo_data(30),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(30),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_29x: FDE port map (
      Q => cpo_data(29),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(29),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_28x: FDE port map (
      Q => cpo_data(28),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(28),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_27x: FDE port map (
      Q => cpo_data(27),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(27),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_26x: FDE port map (
      Q => cpo_data(26),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(26),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_25x: FDE port map (
      Q => cpo_data(25),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(25),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_24x: FDE port map (
      Q => cpo_data(24),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(24),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_23x: FDE port map (
      Q => cpo_data(23),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(23),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_22x: FDE port map (
      Q => cpo_data(22),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(22),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_21x: FDE port map (
      Q => cpo_data(21),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(21),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_20x: FDE port map (
      Q => cpo_data(20),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(20),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_19x: FDE port map (
      Q => cpo_data(19),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(19),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_18x: FDE port map (
      Q => cpo_data(18),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(18),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_17x: FDE port map (
      Q => cpo_data(17),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(17),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_16x: FDE port map (
      Q => cpo_data(16),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(16),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_15x: FDE port map (
      Q => cpo_data(15),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(15),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_14x: FDE port map (
      Q => cpo_data(14),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(14),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_13x: FDE port map (
      Q => cpo_data(13),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(13),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_12x: FDE port map (
      Q => cpo_data(12),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(12),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_11x: FDE port map (
      Q => cpo_data(11),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(11),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_10x: FDE port map (
      Q => cpo_data(10),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(10),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_9x: FDE port map (
      Q => cpo_data(9),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(9),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_8x: FDE port map (
      Q => cpo_data(8),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(8),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_7x: FDE port map (
      Q => cpo_data(7),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(7),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_6x: FDE port map (
      Q => cpo_data(6),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(6),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_5x: FDE port map (
      Q => cpo_data(5),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(5),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_4x: FDE port map (
      Q => cpo_data(4),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(4),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_3x: FDE port map (
      Q => cpo_data(3),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(3),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_2x: FDE port map (
      Q => cpo_data(2),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(2),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_1x: FDE port map (
      Q => cpo_data(1),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(1),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_e_stdata_0x: FDE port map (
      Q => cpo_data(0),
      D => GRLFPC2_0_COMB_V_E_STDATA_1(0),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_fsr_nonstd: FDE port map (
      Q => GRLFPC2_0_R_FSR_NONSTD,
      D => GRLFPC2_0_COMB_V_FSR_NONSTD_1,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_fsr_rd_1x: FDE port map (
      Q => GRLFPC2_0_R_FSR_RD(1),
      D => GRLFPC2_0_COMB_V_FSR_RD_1(1),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_fsr_rd_0x: FDE port map (
      Q => GRLFPC2_0_R_FSR_RD(0),
      D => GRLFPC2_0_COMB_V_FSR_RD_1(0),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_fsr_tem_4x: FDE port map (
      Q => GRLFPC2_0_R_FSR_TEM(4),
      D => GRLFPC2_0_COMB_V_FSR_TEM_1(4),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_fsr_tem_3x: FDE port map (
      Q => GRLFPC2_0_R_FSR_TEM(3),
      D => GRLFPC2_0_COMB_V_FSR_TEM_1(3),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_fsr_tem_2x: FDE port map (
      Q => GRLFPC2_0_R_FSR_TEM(2),
      D => GRLFPC2_0_COMB_V_FSR_TEM_1(2),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_fsr_tem_1x: FDE port map (
      Q => GRLFPC2_0_R_FSR_TEM(1),
      D => GRLFPC2_0_COMB_V_FSR_TEM_1(1),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_fsr_tem_0x: FDE port map (
      Q => GRLFPC2_0_R_FSR_TEM(0),
      D => GRLFPC2_0_COMB_V_FSR_TEM_1(0),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_a_rs1d: FDE port map (
      Q => GRLFPC2_0_R_A_RS1D,
      D => GRLFPC2_0_COMB_RS1D_1,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_a_rs2d: FDE port map (
      Q => GRLFPC2_0_R_A_RS2D,
      D => GRLFPC2_0_N_718_I,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_a_rf2ren_1x: FDE port map (
      Q => GRLFPC2_0_R_A_RF2REN(1),
      D => GRLFPC2_0_N_703,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_a_rf2ren_2x: FDE port map (
      Q => GRLFPC2_0_R_A_RF2REN(2),
      D => GRLFPC2_0_N_657_I,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_fsr_ftt_0x: FDE port map (
      Q => GRLFPC2_0_R_FSR_FTT(0),
      D => GRLFPC2_0_N_721_I,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_fsr_ftt_2x: FDE port map (
      Q => GRLFPC2_0_R_FSR_FTT(2),
      D => GRLFPC2_0_N_720_I,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_a_rf1ren_1x: FDE port map (
      Q => GRLFPC2_0_R_A_RF1REN(1),
      D => GRLFPC2_0_N_637,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_a_rf1ren_2x: FDE port map (
      Q => GRLFPC2_0_R_A_RF1REN(2),
      D => GRLFPC2_0_N_615,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_state_1x: FDE port map (
      Q => GRLFPC2_0_R_STATE(1),
      D => GRLFPC2_0_COMB_V_STATE_1(1),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_state_0x: FDE port map (
      Q => GRLFPC2_0_R_STATE(0),
      D => GRLFPC2_0_COMB_V_STATE_1(0),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_fsr_fcc_1x: FDE port map (
      Q => CPO_CC_1_INT_4,
      D => GRLFPC2_0_COMB_V_FSR_FCC_1(1),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_fsr_fcc_0x: FDE port map (
      Q => CPO_CC_0_INT_3,
      D => GRLFPC2_0_COMB_V_FSR_FCC_1(0),
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_i_exec: FDE port map (
      Q => GRLFPC2_0_R_I_EXEC,
      D => GRLFPC2_0_N_602,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_fsr_aexc_4x: FDE port map (
      Q => GRLFPC2_0_R_FSR_AEXC(4),
      D => GRLFPC2_0_N_728_I,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_fsr_aexc_3x: FDE port map (
      Q => GRLFPC2_0_R_FSR_AEXC(3),
      D => GRLFPC2_0_N_729_I,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_fsr_aexc_2x: FDE port map (
      Q => GRLFPC2_0_R_FSR_AEXC(2),
      D => GRLFPC2_0_N_730_I,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_fsr_aexc_1x: FDE port map (
      Q => GRLFPC2_0_R_FSR_AEXC(1),
      D => GRLFPC2_0_N_731_I,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_fsr_aexc_0x: FDE port map (
      Q => GRLFPC2_0_R_FSR_AEXC(0),
      D => GRLFPC2_0_N_732_I,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_fsr_cexc_4x: FDE port map (
      Q => GRLFPC2_0_R_FSR_CEXC(4),
      D => GRLFPC2_0_N_723_I,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_fsr_cexc_3x: FDE port map (
      Q => GRLFPC2_0_R_FSR_CEXC(3),
      D => GRLFPC2_0_N_724_I,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_fsr_cexc_2x: FDE port map (
      Q => GRLFPC2_0_R_FSR_CEXC(2),
      D => GRLFPC2_0_N_725_I,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_fsr_cexc_1x: FDE port map (
      Q => GRLFPC2_0_R_FSR_CEXC(1),
      D => GRLFPC2_0_N_726_I,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_fsr_cexc_0x: FDE port map (
      Q => GRLFPC2_0_R_FSR_CEXC(0),
      D => GRLFPC2_0_N_727_I,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_a_afq: FDE port map (
      Q => GRLFPC2_0_R_A_AFQ,
      D => GRLFPC2_0_COMB_V_A_AFQ_1,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_a_fpop: FDE port map (
      Q => GRLFPC2_0_R_A_FPOP,
      D => GRLFPC2_0_COMB_FPOP_1,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_a_ld: FDE port map (
      Q => GRLFPC2_0_R_A_LD,
      D => GRLFPC2_0_COMB_V_A_LD_1,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_a_st: FDE port map (
      Q => GRLFPC2_0_R_A_ST,
      D => GRLFPC2_0_COMB_V_A_ST_1,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_r_a_afsr: FDE port map (
      Q => GRLFPC2_0_R_A_AFSR,
      D => GRLFPC2_0_COMB_V_A_AFSR_1,
      C => clk,
      CE => holdn);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_372x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(372),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23(113),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_373x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(373),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_MIXOIN_3_I(0),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_377x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(377),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_NOTREMBIT(3),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_357x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(357),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1766_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_358x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(358),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1765_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_359x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(359),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1764_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_360x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(360),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1763_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_361x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(361),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1762_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_362x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(362),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1761_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_363x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(363),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1760_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_364x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(364),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1759_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_365x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(365),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1758_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_366x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(366),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1757_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_367x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(367),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1756_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_368x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(368),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1755_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_369x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(369),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1754_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_370x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(370),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1753_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_371x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(371),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1752_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_342x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(342),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1781_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_343x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(343),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1780_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_344x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(344),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1779_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_345x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(345),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1778_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_346x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(346),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1777_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_347x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(347),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1776_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_348x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(348),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1775_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_349x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(349),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1774_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_350x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(350),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1773_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_351x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(351),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1772_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_352x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(352),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1771_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_353x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(353),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1770_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_354x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(354),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1769_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_355x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(355),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1768_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_356x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(356),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1767_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_327x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(327),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1796_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_328x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(328),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1795_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_329x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(329),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1794_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_330x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(330),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1793_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_331x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(331),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1792_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_332x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(332),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1791_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_333x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(333),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1790_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_334x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(334),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1789_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_335x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(335),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1788_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_336x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(336),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1787_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_337x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(337),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1786_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_338x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(338),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1785_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_339x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(339),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1784_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_340x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(340),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1783_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_341x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(341),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1782_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_312x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(312),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(53),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_313x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(313),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(54),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_314x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(314),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(55),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_315x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(315),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1724_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_316x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(316),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1751_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_317x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(317),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1806_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_318x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(318),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1805_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_319x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(319),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_23_I_I(60),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_320x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(320),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1803_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_321x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(321),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1802_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_322x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(322),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1801_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_323x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(323),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1800_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_324x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(324),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1799_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_325x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(325),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1798_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_326x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(326),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1797_I,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_297x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(297),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(38),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_298x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(298),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(39),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_299x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(299),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(40),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_300x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(300),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(41),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_301x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(301),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(42),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_302x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(302),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(43),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_303x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(303),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(44),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_304x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(304),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(45),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_305x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(305),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(46),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_306x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(306),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(47),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_307x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(307),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(48),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_308x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(308),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(49),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_309x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(309),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(50),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_310x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(310),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(51),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_311x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(311),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(52),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_282x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(282),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(23),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_283x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(283),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(24),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_284x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(284),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(25),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_285x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(285),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(26),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_286x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(286),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(27),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_287x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(287),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(28),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_288x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(288),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(29),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_289x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(289),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(30),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_290x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(290),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(31),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_291x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(291),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(32),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_292x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(292),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(33),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_293x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(293),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(34),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_294x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(294),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(35),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_295x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(295),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(36),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_296x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(296),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(37),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_267x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(267),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(8),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_268x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(268),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(9),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_269x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(269),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(10),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_270x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(270),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(11),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_271x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(271),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(12),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_272x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(272),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(13),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_273x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(273),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(14),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_274x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(274),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(15),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_275x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(275),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(16),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_276x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(276),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(17),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_277x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(277),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(18),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_278x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(278),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(19),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_279x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(279),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(20),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_280x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(280),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(21),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_281x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(281),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(22),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_252x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(252),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(252),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_253x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(253),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(253),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_254x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(254),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(254),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_255x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(255),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(255),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_256x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(256),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(256),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_257x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(257),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(257),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_258x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(258),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_49(258),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_259x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(259),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(0),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_260x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(260),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(1),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_261x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(261),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(2),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_262x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(262),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(3),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_263x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(263),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(4),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_264x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(264),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(5),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_265x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(265),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(6),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_266x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(266),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_DPATH_NEW_8(7),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_UN2_NOTABORTWB_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_237x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(237),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(237),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_238x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(238),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(238),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_239x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(239),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(239),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_240x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(240),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(240),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_241x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(241),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(241),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_242x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(242),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(242),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_243x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(243),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(243),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_244x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(244),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(244),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_247x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(247),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(247),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_248x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(248),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(248),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_249x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(249),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(249),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_250x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(250),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(250),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_251x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(251),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(251),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_222x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(222),
      D => GRLFPC2_0_FPO_FRAC(9),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_223x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(223),
      D => GRLFPC2_0_FPO_FRAC(8),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_224x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(224),
      D => GRLFPC2_0_FPO_FRAC(7),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_225x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(225),
      D => GRLFPC2_0_FPO_FRAC(6),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_226x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(226),
      D => GRLFPC2_0_FPO_FRAC(5),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_227x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(227),
      D => GRLFPC2_0_FPO_FRAC(4),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_228x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(228),
      D => GRLFPC2_0_FPO_FRAC(3),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_229x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(229),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_225,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_230x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(230),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_224,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_231x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(231),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_223,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_207x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(207),
      D => GRLFPC2_0_FPO_FRAC(24),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_208x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(208),
      D => GRLFPC2_0_FPO_FRAC(23),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_209x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(209),
      D => GRLFPC2_0_FPO_FRAC(22),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_210x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(210),
      D => GRLFPC2_0_FPO_FRAC(21),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_211x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(211),
      D => GRLFPC2_0_FPO_FRAC(20),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_212x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(212),
      D => GRLFPC2_0_FPO_FRAC(19),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_213x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(213),
      D => GRLFPC2_0_FPO_FRAC(18),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_214x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(214),
      D => GRLFPC2_0_FPO_FRAC(17),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_215x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(215),
      D => GRLFPC2_0_FPO_FRAC(16),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_216x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(216),
      D => GRLFPC2_0_FPO_FRAC(15),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_217x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(217),
      D => GRLFPC2_0_FPO_FRAC(14),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_218x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(218),
      D => GRLFPC2_0_FPO_FRAC(13),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_219x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(219),
      D => GRLFPC2_0_FPO_FRAC(12),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_220x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(220),
      D => GRLFPC2_0_FPO_FRAC(11),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_221x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(221),
      D => GRLFPC2_0_FPO_FRAC(10),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_192x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(192),
      D => GRLFPC2_0_FPO_FRAC(39),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_193x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(193),
      D => GRLFPC2_0_FPO_FRAC(38),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_194x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(194),
      D => GRLFPC2_0_FPO_FRAC(37),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_195x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(195),
      D => GRLFPC2_0_FPO_FRAC(36),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_196x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(196),
      D => GRLFPC2_0_FPO_FRAC(35),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_197x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(197),
      D => GRLFPC2_0_FPO_FRAC(34),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_198x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(198),
      D => GRLFPC2_0_FPO_FRAC(33),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_199x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(199),
      D => GRLFPC2_0_FPO_FRAC(32),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_200x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(200),
      D => GRLFPC2_0_FPO_FRAC(31),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_201x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(201),
      D => GRLFPC2_0_FPO_FRAC(30),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_202x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(202),
      D => GRLFPC2_0_FPO_FRAC(29),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_203x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(203),
      D => GRLFPC2_0_FPO_FRAC(28),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_204x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(204),
      D => GRLFPC2_0_FPO_FRAC(27),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_205x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(205),
      D => GRLFPC2_0_FPO_FRAC(26),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_206x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(206),
      D => GRLFPC2_0_FPO_FRAC(25),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_177x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(177),
      D => GRLFPC2_0_FPO_FRAC(54),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_178x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(178),
      D => GRLFPC2_0_FPO_FRAC(53),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_179x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(179),
      D => GRLFPC2_0_FPO_FRAC(52),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_180x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(180),
      D => GRLFPC2_0_FPO_FRAC(51),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_181x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(181),
      D => GRLFPC2_0_FPO_FRAC(50),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_182x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(182),
      D => GRLFPC2_0_FPO_FRAC(49),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_183x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(183),
      D => GRLFPC2_0_FPO_FRAC(48),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_184x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(184),
      D => GRLFPC2_0_FPO_FRAC(47),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_185x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(185),
      D => GRLFPC2_0_FPO_FRAC(46),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_186x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(186),
      D => GRLFPC2_0_FPO_FRAC(45),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_187x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(187),
      D => GRLFPC2_0_FPO_FRAC(44),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_188x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(188),
      D => GRLFPC2_0_FPO_FRAC(43),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_189x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(189),
      D => GRLFPC2_0_FPO_FRAC(42),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_190x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(190),
      D => GRLFPC2_0_FPO_FRAC(41),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_191x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(191),
      D => GRLFPC2_0_FPO_FRAC(40),
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_174x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(174),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2276,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_175x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(175),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_279,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_176x: FDE port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(176),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_278,
      C => clk,
      CE => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_XZTREGLOADEN);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_102x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(102),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(102),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_103x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(103),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(103),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_104x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(104),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(104),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_105x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(105),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(105),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_106x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(106),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(106),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_107x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(107),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(107),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_108x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(108),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(108),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_109x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(109),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(109),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_110x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(110),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(110),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_111x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(111),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(111),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_112x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(112),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(112),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_113x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(113),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(113),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_114x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(114),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(114),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_87x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(87),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(87),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_88x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(88),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(88),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_89x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(89),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(89),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_90x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(90),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(90),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_91x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(91),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(91),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_92x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(92),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(92),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_93x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(93),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(93),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_94x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(94),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(94),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_95x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(95),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(95),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_96x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(96),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(96),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_97x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(97),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(97),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_98x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(98),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(98),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_99x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(99),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(99),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_100x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(100),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(100),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_101x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(101),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(101),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_72x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(72),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(72),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_73x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(73),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(73),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_74x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(74),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(74),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_75x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(75),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_76x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(76),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_77x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(77),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(77),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_78x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(78),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(78),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_79x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(79),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(79),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_80x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(80),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(80),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_81x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(81),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(81),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_82x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(82),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(82),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_83x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(83),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_84x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(84),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(84),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_85x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(85),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(85),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_86x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(86),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(86),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_58x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(58),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(58),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_59x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(59),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(59),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_60x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(60),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(60),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_61x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(61),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(61),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_62x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(62),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(62),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_63x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(63),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(63),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_64x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(64),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_65x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(65),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(65),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_66x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(66),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_67x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(67),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(67),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_68x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(68),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(68),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_69x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(69),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(69),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_70x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(70),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(70),
      C => clk);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpath_71x: FD port map (
      Q => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(71),
      D => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_RIN_DPATH(71),
      C => clk);
  x_I_768: INV port map (
      I => rst,
      O => RST_I);
  x_I_767: INV port map (
      I => cpi_d_inst(31),
      O => CPI_D_INST_I(31));
  x_I_766: INV port map (
      I => holdn,
      O => HOLDN_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_cry_55_ma: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(55),
      I1 => NN_2,
      LO => N_20279);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_cry_55_ma: MULT_AND port map (
      I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(55),
      I1 => NN_2,
      LO => N_20281);
  x_grlfpc2_0_comb_v_fsr_N_727_i: LUT4_L 
  generic map(
    INIT => X"F777"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_FSR_N_727_I_1,
    I1 => GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_0(0),
    I2 => GRLFPC2_0_R_FSR_CEXC(0),
    I3 => GRLFPC2_0_V_FSR_CEXC_3_SQMUXA,
    LO => GRLFPC2_0_N_727_I);
  x_grlfpc2_0_comb_v_fsr_N_726_i: LUT4_L 
  generic map(
    INIT => X"F777"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_FSR_N_726_I_1,
    I1 => GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_0(1),
    I2 => GRLFPC2_0_R_FSR_CEXC(1),
    I3 => GRLFPC2_0_V_FSR_CEXC_3_SQMUXA,
    LO => GRLFPC2_0_N_726_I);
  x_grlfpc2_0_comb_v_fsr_N_725_i: LUT4_L 
  generic map(
    INIT => X"F777"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_FSR_N_725_I_1,
    I1 => GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_0(2),
    I2 => GRLFPC2_0_R_FSR_CEXC(2),
    I3 => GRLFPC2_0_V_FSR_CEXC_3_SQMUXA,
    LO => GRLFPC2_0_N_725_I);
  x_grlfpc2_0_comb_v_fsr_N_724_i: LUT4_L 
  generic map(
    INIT => X"F777"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_FSR_N_724_I_1,
    I1 => GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_0(3),
    I2 => GRLFPC2_0_R_FSR_CEXC(3),
    I3 => GRLFPC2_0_V_FSR_CEXC_3_SQMUXA,
    LO => GRLFPC2_0_N_724_I);
  x_grlfpc2_0_comb_v_fsr_N_723_i: LUT4_L 
  generic map(
    INIT => X"F777"
  )
  port map (
    I0 => GRLFPC2_0_COMB_V_FSR_N_723_I_1,
    I1 => GRLFPC2_0_COMB_V_FSR_CEXC_1_IV_0(4),
    I2 => GRLFPC2_0_R_FSR_CEXC(4),
    I3 => GRLFPC2_0_V_FSR_CEXC_3_SQMUXA,
    LO => GRLFPC2_0_N_723_I);
  x_grlfpc2_0_comb_v_x_ld_1: LUT3_L 
  generic map(
    INIT => X"02"
  )
  port map (
    I0 => GRLFPC2_0_R_M_LD,
    I1 => cpi_m_trap,
    I2 => cpi_m_annul,
    LO => GRLFPC2_0_COMB_V_X_LD_1);
  x_grlfpc2_0_comb_v_x_fpop_1: LUT3_L 
  generic map(
    INIT => X"02"
  )
  port map (
    I0 => GRLFPC2_0_R_M_FPOP,
    I1 => cpi_m_trap,
    I2 => cpi_m_annul,
    LO => GRLFPC2_0_COMB_V_X_FPOP_1);
  x_grlfpc2_0_comb_v_x_afsr_1: LUT3_L 
  generic map(
    INIT => X"02"
  )
  port map (
    I0 => GRLFPC2_0_R_M_AFSR,
    I1 => cpi_m_trap,
    I2 => cpi_m_annul,
    LO => GRLFPC2_0_COMB_V_X_AFSR_1);
  x_grlfpc2_0_comb_v_x_afq_1: LUT3_L 
  generic map(
    INIT => X"02"
  )
  port map (
    I0 => GRLFPC2_0_R_M_AFQ,
    I1 => cpi_m_trap,
    I2 => cpi_m_annul,
    LO => GRLFPC2_0_COMB_V_X_AFQ_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_m_0_4_rep1: LUT4_L 
  generic map(
    INIT => X"7545"
  )
  port map (
    I0 => N_13323,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(4),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_4_REP1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_m_0_7_rep1: LUT4_L 
  generic map(
    INIT => X"40FB"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(7),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_M_0_1(7),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_7_REP1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_m_0_2_rep1: LUT4_L 
  generic map(
    INIT => X"40FB"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(2),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_M_0_1(2),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_2_REP1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_m_0_3_rep1: LUT4_L 
  generic map(
    INIT => X"25EA"
  )
  port map (
    I0 => N_12615,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_371,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_M_0_1(3),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_3_REP1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_m_0_5_rep1: LUT4_L 
  generic map(
    INIT => X"40FB"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(5),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_M_0_1(5),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_5_REP1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_m_0_6_rep1: LUT4_L 
  generic map(
    INIT => X"40FB"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(6),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_M_0_1(6),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_6_REP1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_m_0_0_rep1: LUT4_L 
  generic map(
    INIT => X"40FB"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(0),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_M_0_1(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_0_REP1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_m_0_1_rep1: LUT4_L 
  generic map(
    INIT => X"40FB"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_M_0_1(1),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_1_REP1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_1_i: LUT4_L 
  generic map(
    INIT => X"DFFF"
  )
  port map (
    I0 => N_15852,
    I1 => N_15853,
    I2 => N_15854,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_1_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_1_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_2_i: LUT4_L 
  generic map(
    INIT => X"DFFF"
  )
  port map (
    I0 => N_15820,
    I1 => N_15821,
    I2 => N_15822,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_2_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_2_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_3_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => N_15883,
    I1 => N_15884,
    I2 => N_15885,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_3_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_3_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_4_i: LUT4_L 
  generic map(
    INIT => X"DFFF"
  )
  port map (
    I0 => N_15896,
    I1 => N_15897,
    I2 => N_15898,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_4_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_4_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_5_i: LUT4_L 
  generic map(
    INIT => X"FF7F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_5_I_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_5_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_5_3,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M_0(51),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_5_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_6_i: LUT4_L 
  generic map(
    INIT => X"EFFF"
  )
  port map (
    I0 => N_13133,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_NOTSRRES_M(53),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_6_I_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_6_2,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_6_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_7_i: LUT4_L 
  generic map(
    INIT => X"DFFF"
  )
  port map (
    I0 => N_15807,
    I1 => N_15808,
    I2 => N_15809,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_7_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_7_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_8_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => N_15775,
    I1 => N_15776,
    I2 => N_15777,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_8_2,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_8_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_9_i: LUT4_L 
  generic map(
    INIT => X"FFBF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_9_I_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_9_2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_9_6_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M_0(56),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_9_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_21_i: LUT4_L 
  generic map(
    INIT => X"FF7F"
  )
  port map (
    I0 => N_12973,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_21_I_1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_21_3,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M(42),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_21_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_22_i: LUT4_L 
  generic map(
    INIT => X"75FF"
  )
  port map (
    I0 => N_13217,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(43),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_22_5,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_22_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_23_i: LUT4_L 
  generic map(
    INIT => X"FF7F"
  )
  port map (
    I0 => N_13005,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_23_I_1_0,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_23_3,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2_M(44),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_23_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_24_i: LUT4_L 
  generic map(
    INIT => X"75FF"
  )
  port map (
    I0 => N_13154,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(45),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_24_5,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_24_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_30_i: LUT4_L 
  generic map(
    INIT => X"BFFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_30_I_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_30_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_30_4,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_30_7,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_30_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_40_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_40_I_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_40_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_40_2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_40_5,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_40_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_47_i: LUT4_L 
  generic map(
    INIT => X"7FFF"
  )
  port map (
    I0 => N_13061,
    I1 => N_15367,
    I2 => N_15368,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_47_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_47_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_48_i: LUT4_L 
  generic map(
    INIT => X"75FF"
  )
  port map (
    I0 => N_13175,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(9),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_48_5,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_48_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_51_i: LUT4_L 
  generic map(
    INIT => X"BFFF"
  )
  port map (
    I0 => N_13086,
    I1 => N_13088,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_51_I_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_51_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_51_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_52_i: LUT4_L 
  generic map(
    INIT => X"75FF"
  )
  port map (
    I0 => N_13196,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(13),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_52_5,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_52_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_53_i: LUT4_L 
  generic map(
    INIT => X"BFFF"
  )
  port map (
    I0 => N_13111,
    I1 => N_13113,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_53_I_1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_53_3,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_53_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_54_i: LUT4_L 
  generic map(
    INIT => X"75FF"
  )
  port map (
    I0 => N_13238,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_S_2(15),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_54_5,
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_54_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r_dpaths_55_i: LUT4_L 
  generic map(
    INIT => X"BF3F"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_DPATH_NEW_8_SQMUXA,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_55_I_1,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHSR_55_2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_S_1_2(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATHS_55_I);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_m_0_0x: LUT4_L 
  generic map(
    INIT => X"40FB"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(0),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_M_0_1(0),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT(0));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_m_0_1x: LUT4_L 
  generic map(
    INIT => X"40FB"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(1),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_M_0_1(1),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT(1));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_m_0_2x: LUT4_L 
  generic map(
    INIT => X"40FB"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(2),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_M_0_1(2),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT(2));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_m_0_3x: LUT4_L 
  generic map(
    INIT => X"25EA"
  )
  port map (
    I0 => N_12615,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_371,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_M_0_1(3),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT(3));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_m_0_4x: LUT4_L 
  generic map(
    INIT => X"7545"
  )
  port map (
    I0 => N_13323,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_3,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(4),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT(4));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_m_0_5x: LUT4_L 
  generic map(
    INIT => X"40FB"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(5),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_M_0_1(5),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT(5));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_m_0_6x: LUT4_L 
  generic map(
    INIT => X"40FB"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(6),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_M_0_1(6),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT(6));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_pxs_multiplexormulxff_result_m_0_7x: LUT4_L 
  generic map(
    INIT => X"40FB"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_RN_3,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_NOTSQRTLFTCC_1_28_0_SN,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT1(7),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT_M_0_1(7),
    LO => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_PXS_MULTIPLEXORMULXFF_RESULT(7));
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_56: LUT4 
  generic map(
    INIT => X"8778"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(59),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(56),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_56);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_55: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(55),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(55),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_55);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_54: LUT4 
  generic map(
    INIT => X"8778"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(61),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(54),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_54);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_53: LUT4 
  generic map(
    INIT => X"8778"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(62),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(53),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_53);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_52: LUT4 
  generic map(
    INIT => X"8778"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(63),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(52),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_52);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_51: LUT4 
  generic map(
    INIT => X"8778"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(51),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_51);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_50: LUT4 
  generic map(
    INIT => X"8778"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(65),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(50),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_50);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_49: LUT4 
  generic map(
    INIT => X"8778"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(49),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_49);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_48: LUT4 
  generic map(
    INIT => X"8778"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(67),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(48),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_48);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_47: LUT4 
  generic map(
    INIT => X"8778"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(68),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(47),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_47);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_46: LUT4 
  generic map(
    INIT => X"8778"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(69),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(46),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_46);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_45: LUT4 
  generic map(
    INIT => X"8778"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(70),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(45),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_45);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_44: LUT4 
  generic map(
    INIT => X"8778"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(71),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(44),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_44);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_43: LUT4 
  generic map(
    INIT => X"8778"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(72),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(43),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_43);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_42: LUT4 
  generic map(
    INIT => X"8778"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(73),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(42),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_42);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_41: LUT4 
  generic map(
    INIT => X"8778"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(74),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(41),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_41);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_40: LUT4 
  generic map(
    INIT => X"8778"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(40),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_40);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_39: LUT4 
  generic map(
    INIT => X"8778"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(39),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_39);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_38: LUT4 
  generic map(
    INIT => X"8778"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(77),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(38),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_38);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_37: LUT4 
  generic map(
    INIT => X"8778"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(78),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(37),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_37);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_36: LUT4 
  generic map(
    INIT => X"8778"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(79),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(36),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_36);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_35: LUT4 
  generic map(
    INIT => X"8778"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(80),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(35),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_35);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_34: LUT4 
  generic map(
    INIT => X"8778"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(81),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(34),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_34);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_33: LUT4 
  generic map(
    INIT => X"8778"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(82),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(33),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_33);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_32: LUT4 
  generic map(
    INIT => X"8778"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(32),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ_I(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_32);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_31: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(31),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(31),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_31);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_30: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_30);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_29: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(29),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(29),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_29);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_28: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(28),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(28),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_28);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_27: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(27),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(27),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_27);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_26: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(26),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(26),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_26);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_25: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(25),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(25),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_25);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_24: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(24),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(24),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_24);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_23: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(23),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(23),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_23);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_22: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(22),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(22),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_22);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_21: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(21),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(21),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_21);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_20: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(20),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(20),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_20);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_19: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(19),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(19),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_19);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_18: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(18),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(18),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_18);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_17: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(17),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_17);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_16: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(16),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(16),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_16);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_15: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(15),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(15),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_15);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_14: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(14),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(14),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_14);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_13: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(13),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(13),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_13);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_12: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(12),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(12),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_12);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_11: LUT4 
  generic map(
    INIT => X"B847"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_118,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(46),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_11_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_11);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_10: LUT4 
  generic map(
    INIT => X"B847"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_117,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(47),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_10_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_10);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_9: LUT4 
  generic map(
    INIT => X"B847"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_116,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(48),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_9_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_9);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_8: LUT4 
  generic map(
    INIT => X"B847"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_115,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(49),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_8_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_8);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_7: LUT4 
  generic map(
    INIT => X"B847"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_114,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(50),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_7_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_6: LUT4 
  generic map(
    INIT => X"B847"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_113,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(51),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_6_1,
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_5: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(5),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_4: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(4),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_3: LUT3 
  generic map(
    INIT => X"69"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_C_FAX_XZYBUS(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_2: LUT4 
  generic map(
    INIT => X"9A95"
  )
  port map (
    I0 => N_13011,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_109,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_2261_I,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(55),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_1: LUT2 
  generic map(
    INIT => X"6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN20_XZXBUS(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r1_un6_grfpuf_axb_0: LUT4 
  generic map(
    INIT => X"639C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN39_XZYBUSLSBS,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_2_1(0),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R1_UN6_GRFPUF_AXB_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_56: LUT3 
  generic map(
    INIT => X"87"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(59),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_56);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_55: LUT4 
  generic map(
    INIT => X"B847"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(60),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(18),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_55);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_54: LUT3 
  generic map(
    INIT => X"87"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(61),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_54);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_53: LUT3 
  generic map(
    INIT => X"87"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(62),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_53);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_52: LUT3 
  generic map(
    INIT => X"87"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(63),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_52);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_51: LUT3 
  generic map(
    INIT => X"87"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(64),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_51);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_50: LUT3 
  generic map(
    INIT => X"87"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(65),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_50);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_49: LUT3 
  generic map(
    INIT => X"87"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(66),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_49);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_48: LUT3 
  generic map(
    INIT => X"87"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(67),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_48);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_47: LUT3 
  generic map(
    INIT => X"87"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(68),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_47);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_46: LUT3 
  generic map(
    INIT => X"87"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(69),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_46);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_45: LUT3 
  generic map(
    INIT => X"87"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(70),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(17),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_45);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_44: LUT3 
  generic map(
    INIT => X"87"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(71),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_44);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_43: LUT3 
  generic map(
    INIT => X"87"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(72),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_43);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_42: LUT3 
  generic map(
    INIT => X"87"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(73),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_42);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_41: LUT3 
  generic map(
    INIT => X"87"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(74),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_41);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_40: LUT3 
  generic map(
    INIT => X"87"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(75),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_40);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_39: LUT3 
  generic map(
    INIT => X"87"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(76),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_39);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_38: LUT3 
  generic map(
    INIT => X"87"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(77),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_38);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_37: LUT3 
  generic map(
    INIT => X"87"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(78),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_37);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_36: LUT3 
  generic map(
    INIT => X"87"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(79),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_36);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_35: LUT3 
  generic map(
    INIT => X"87"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(80),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_35);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_34: LUT3 
  generic map(
    INIT => X"87"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(81),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_34);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_33: LUT3 
  generic map(
    INIT => X"87"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(82),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_33);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_32: LUT3 
  generic map(
    INIT => X"87"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(83),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_32);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_31: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(31),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_31);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_30: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(85),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_30);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_29: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(86),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_29);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_28: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(87),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_28);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_27: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(88),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_27);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_26: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(89),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_26);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_25: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(90),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_25);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_24: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(91),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_24);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_23: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(92),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_23);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_22: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(93),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_22);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_21: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(94),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_21);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_20: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(95),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_20);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_19: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(96),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_19);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_18: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(97),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_18);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_17: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(98),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP2,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_17);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_16: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(99),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_16);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_15: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(100),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_15);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_14: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(101),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_14);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_13: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(102),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_13);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_12: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(103),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_12);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_11: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(104),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_11);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_10: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(105),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_10);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_9: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(106),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_9);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_8: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(107),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_8);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_7: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(108),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_6: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(109),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_5: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(110),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_4: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(111),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_3: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(30),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(112),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_2: LUT4 
  generic map(
    INIT => X"CA35"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS_2(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(113),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL_17_REP1,
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_1: LUT2 
  generic map(
    INIT => X"6"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN20_XZXBUS(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(1),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_r0_un6_grfpuf_axb_0: LUT4 
  generic map(
    INIT => X"639C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_UN39_XZYBUSLSBS,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZXBUS(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_FAX_XZYBUS_2_1(0),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_WAITQ(0),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R0_UN6_GRFPUF_AXB_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_axb_11: LUT4 
  generic map(
    INIT => X"936C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_999,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_1(11),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_11);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_axb_10: LUT4 
  generic map(
    INIT => X"936C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_998,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_1(10),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(33),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_10);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_axb_9: LUT4 
  generic map(
    INIT => X"936C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1021,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(9),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_9);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_axb_8: LUT4 
  generic map(
    INIT => X"936C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1020,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(8),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_8);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_axb_7: LUT4 
  generic map(
    INIT => X"936C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1019,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(7),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_axb_6: LUT3 
  generic map(
    INIT => X"96"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(6),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_1(6),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_axb_5: LUT4 
  generic map(
    INIT => X"936C"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_N_1017,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(5),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(31),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_axb_4: LUT3 
  generic map(
    INIT => X"96"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(4),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_EXPYBUS_1(4),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_axb_3: LUT3 
  generic map(
    INIT => X"96"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(3),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(3),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_axb_2: LUT3 
  generic map(
    INIT => X"96"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(2),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(2),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_axb_1: LUT3 
  generic map(
    INIT => X"96"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(1),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un6_grfpue_axb_0: LUT3 
  generic map(
    INIT => X"96"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_DPXX_LEFTSHIFTERBL_SLCONTROL(0),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_EXPADDERSHFT_EXPXBUS(0),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN6_GRFPUE_AXB_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_axb_6: LUT1 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(79),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_axb_5: LUT1 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(80),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_axb_4: LUT1 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(81),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_axb_3: LUT1 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(82),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_axb_2: LUT1 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(83),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_axb_1: LUT1 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(84),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_un1_notsampledwait_axb_0: LUT1 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_PCTRL(85),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_UN1_NOTSAMPLEDWAIT_AXB_0);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_axb_11: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(233),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(246),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_11);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_axb_10: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(234),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(247),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_10);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_axb_9: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(235),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(248),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_9);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_axb_8: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(236),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(249),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_8);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_axb_7: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(237),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(250),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_7);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_axb_6: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(238),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(251),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_6);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_axb_5: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(239),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(252),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_5);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_axb_4: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(240),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(253),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_4);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_axb_3: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(241),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(254),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_3);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_axb_2: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(242),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(255),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_2);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_grfpue_axb_1: LUT2 
  generic map(
    INIT => X"9"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(243),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(256),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_GRFPUE_AXB_1);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_7_and: LUT3 
  generic map(
    INIT => X"2A"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_7_AND1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(1),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(25),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_7_AND);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_6_and: LUT2 
  generic map(
    INIT => X"2"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_6_AND_1,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(49),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_6_AND);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_5_and: LUT4 
  generic map(
    INIT => X"0001"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(45),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(46),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(47),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(48),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_5_AND);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_4_and: LUT4 
  generic map(
    INIT => X"0001"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(41),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(42),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(43),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(44),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_4_AND);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_3_and: LUT4 
  generic map(
    INIT => X"0001"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(37),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(38),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(39),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(40),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_3_AND);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_2_and: LUT4 
  generic map(
    INIT => X"0001"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(33),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(34),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(35),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(36),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_2_AND);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_1_and: LUT4 
  generic map(
    INIT => X"0001"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(29),
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(30),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(31),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(32),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_1_AND);
  x_grlfpc2_0_grfpul_gen0_grfpulite0_c_inexactsig_un15_inexact_0_and: LUT4 
  generic map(
    INIT => X"0002"
  )
  port map (
    I0 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_NOTAM2_0,
    I1 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(26),
    I2 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(27),
    I3 => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_R_DPATH(28),
    O => GRLFPC2_0_GRFPUL_GEN0_GRFPULITE0_C_INEXACTSIG_UN15_INEXACT_0_AND);
  x_GND: GND port map (
      G => NN_1);
  x_VCC: VCC port map (
      P => NN_2);
  cpo_exc <= CPO_EXC_INT_2;
  cpo_cc(0) <= CPO_CC_0_INT_3;
  cpo_cc(1) <= CPO_CC_1_INT_4;
  rfi1_rd1addr(0) <= RFI2_RD1ADDR_0_INT_5_INT_17;
  rfi1_rd1addr(1) <= RFI2_RD1ADDR_1_INT_6_INT_18;
  rfi1_rd1addr(2) <= RFI2_RD1ADDR_2_INT_7_INT_19;
  rfi1_rd1addr(3) <= RFI2_RD1ADDR_3_INT_8_INT_20;
  rfi1_rd2addr(0) <= RFI2_RD2ADDR_0_INT_9_INT_21;
  rfi1_rd2addr(1) <= RFI2_RD2ADDR_1_INT_10_INT_22;
  rfi1_rd2addr(2) <= RFI2_RD2ADDR_2_INT_11_INT_23;
  rfi1_rd2addr(3) <= RFI2_RD2ADDR_3_INT_12_INT_24;
  rfi1_wraddr(0) <= RFI2_WRADDR_0_INT_13_INT_25;
  rfi1_wraddr(1) <= RFI2_WRADDR_1_INT_14_INT_26;
  rfi1_wraddr(2) <= RFI2_WRADDR_2_INT_15_INT_27;
  rfi1_wraddr(3) <= RFI2_WRADDR_3_INT_16_INT_28;
  rfi2_rd1addr(0) <= RFI2_RD1ADDR_0_INT_5_INT_17;
  rfi2_rd1addr(1) <= RFI2_RD1ADDR_1_INT_6_INT_18;
  rfi2_rd1addr(2) <= RFI2_RD1ADDR_2_INT_7_INT_19;
  rfi2_rd1addr(3) <= RFI2_RD1ADDR_3_INT_8_INT_20;
  rfi2_rd2addr(0) <= RFI2_RD2ADDR_0_INT_9_INT_21;
  rfi2_rd2addr(1) <= RFI2_RD2ADDR_1_INT_10_INT_22;
  rfi2_rd2addr(2) <= RFI2_RD2ADDR_2_INT_11_INT_23;
  rfi2_rd2addr(3) <= RFI2_RD2ADDR_3_INT_12_INT_24;
  rfi2_wraddr(0) <= RFI2_WRADDR_0_INT_13_INT_25;
  rfi2_wraddr(1) <= RFI2_WRADDR_1_INT_14_INT_26;
  rfi2_wraddr(2) <= RFI2_WRADDR_2_INT_15_INT_27;
  rfi2_wraddr(3) <= RFI2_WRADDR_3_INT_16_INT_28;
end beh;

